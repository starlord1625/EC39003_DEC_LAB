CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
380 70 2 80 9
0 76 1536 869
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 76 1536 869
143654930 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 1141 710 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
14 Logic Display~
6 1795 175 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 1821 176 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 1846 175 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 1896 174 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 1871 175 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
7 Ground~
168 1713 636 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
6 74LS83
105 1432 863 0 14 29
0 21 20 19 18 10 11 12 13 2
3 4 5 6 7
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
3 U11
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3747 0 0
0
0
7 Buffer~
58 980 788 0 2 22
0 9 8
0
0 0 624 270
4 4050
-14 -19 14 -11
4 U12A
14 -5 42 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 5 0
1 U
3549 0 0
0
0
7 74LS273
150 1207 750 0 18 37
0 22 8 10 11 12 13 14 15 16
17 21 20 19 18 10 11 12 13
0
0 0 13040 0
7 74LS273
-24 -60 25 -52
3 U10
-11 -61 10 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
10 Ascii Key~
169 1033 162 0 11 12
0 17 16 15 14 52 53 54 9 0
0 57
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
9325 0 0
0
0
7 Ground~
168 1357 840 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
8 3-In OR~
219 1391 538 0 4 22
0 7 24 23 25
0
0 0 624 90
4 4075
-14 -24 14 -16
3 U8A
28 -3 49 5
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
3834 0 0
0
0
9 2-In AND~
219 1416 597 0 3 22
0 5 3 23
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U6D
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 -170575095
65 0 0 0 4 4 3 0
1 U
3363 0 0
0
0
9 2-In AND~
219 1374 599 0 3 22
0 4 3 24
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U6C
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 -120243452
65 0 0 0 4 3 3 0
1 U
7668 0 0
0
0
7 Ground~
168 1543 526 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
6 74LS83
105 1701 555 0 14 29
0 3 4 5 6 2 55 56 2 2
29 28 27 26 57
0
0 0 13040 90
7 74LS83A
-24 -60 25 -52
2 U9
57 -3 71 5
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
7 Ground~
168 1262 379 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
7 74LS157
122 1597 466 0 14 29
0 25 26 6 27 5 28 4 29 3
2 33 32 31 30
0
0 0 13040 602
7 74LS157
-24 -60 25 -52
2 U7
54 -6 68 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3789 0 0
0
0
2 +V
167 1600 59 0 1 3
0 34
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4871 0 0
0
0
9 CA 7-Seg~
184 1600 169 0 18 19
10 36 37 38 39 40 41 42 58 35
0 0 0 0 0 0 0 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3750 0 0
0
0
6 74LS47
187 1573 304 0 14 29
0 30 31 32 33 59 60 42 41 40
39 38 37 36 61
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8778 0 0
0
0
6 74LS47
187 1225 300 0 14 29
0 2 2 2 25 62 63 51 50 49
48 47 46 45 64
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U2
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
538 0 0
0
0
9 CA 7-Seg~
184 1252 165 0 18 19
10 45 46 47 48 49 50 51 65 44
2 0 0 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6843 0 0
0
0
2 +V
167 1252 55 0 1 3
0 43
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3136 0 0
0
0
9 Resistor~
219 1600 109 0 4 5
0 35 34 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
9 Resistor~
219 1252 105 0 4 5
0 44 43 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5670 0 0
0
0
75
0 1 3 0 0 8320 0 0 3 54 0 3
1551 899
1821 899
1821 194
0 1 4 0 0 8320 0 0 4 55 0 3
1541 912
1846 912
1846 193
0 1 5 0 0 8320 0 0 6 56 0 3
1534 929
1871 929
1871 193
0 1 6 0 0 8320 0 0 5 57 0 3
1526 945
1896 945
1896 192
0 1 7 0 0 8320 0 0 2 29 0 3
1517 973
1795 973
1795 193
9 0 2 0 0 4096 0 17 0 0 7 3
1744 589
1744 622
1726 622
8 0 2 0 0 0 0 17 0 0 8 3
1726 589
1726 622
1713 622
5 1 2 0 0 0 0 17 7 0 0 4
1699 589
1699 622
1713 622
1713 630
2 2 8 0 0 8320 0 9 10 0 0 5
980 803
980 837
1124 837
1124 723
1175 723
8 1 9 0 0 4224 0 11 9 0 0 4
1012 186
1012 768
980 768
980 773
0 3 10 0 0 8192 0 0 10 23 0 5
1283 768
1283 846
1138 846
1138 732
1175 732
0 4 11 0 0 8192 0 0 10 22 0 5
1274 777
1274 833
1149 833
1149 741
1175 741
0 5 12 0 0 8192 0 0 10 21 0 5
1262 786
1262 821
1156 821
1156 750
1175 750
0 6 13 0 0 8192 0 0 10 20 0 5
1251 795
1251 812
1167 812
1167 759
1175 759
4 7 14 0 0 4224 0 11 10 0 0 3
1036 186
1036 768
1175 768
3 8 15 0 0 4224 0 11 10 0 0 3
1042 186
1042 777
1175 777
2 9 16 0 0 4224 0 11 10 0 0 3
1048 186
1048 786
1175 786
1 10 17 0 0 4224 0 11 10 0 0 3
1054 186
1054 795
1175 795
9 1 2 0 0 0 0 8 12 0 0 4
1389 833
1389 805
1357 805
1357 834
18 8 13 0 0 4224 0 10 8 0 0 3
1239 795
1407 795
1407 833
17 7 12 0 0 4224 0 10 8 0 0 3
1239 786
1416 786
1416 833
16 6 11 0 0 4224 0 10 8 0 0 3
1239 777
1425 777
1425 833
15 5 10 0 0 4224 0 10 8 0 0 3
1239 768
1434 768
1434 833
14 4 18 0 0 4224 0 10 8 0 0 3
1239 759
1443 759
1443 833
13 3 19 0 0 4224 0 10 8 0 0 3
1239 750
1452 750
1452 833
12 2 20 0 0 4224 0 10 8 0 0 3
1239 741
1461 741
1461 833
11 1 21 0 0 4224 0 10 8 0 0 3
1239 732
1470 732
1470 833
1 1 22 0 0 4224 0 1 10 0 0 3
1153 710
1169 710
1169 714
14 1 7 0 0 128 0 8 13 0 0 8
1389 897
1389 973
1517 973
1517 719
1338 719
1338 567
1385 567
1385 554
3 3 23 0 0 4224 0 13 14 0 0 3
1403 554
1403 573
1415 573
3 2 24 0 0 8320 0 15 13 0 0 3
1373 575
1394 575
1394 553
1 0 4 0 0 0 0 15 0 0 55 3
1364 620
1364 649
1414 649
1 0 5 0 0 0 0 14 0 0 56 3
1406 618
1408 618
1408 635
2 0 3 0 0 0 0 14 0 0 35 3
1424 618
1423 618
1423 656
2 0 3 0 0 0 0 15 0 0 54 3
1382 620
1382 656
1423 656
10 1 2 0 0 0 0 19 16 0 0 4
1551 503
1551 514
1543 514
1543 520
4 0 25 0 0 8320 0 23 0 0 53 4
1239 337
1239 459
1417 459
1417 508
2 13 26 0 0 8320 0 19 17 0 0 4
1623 497
1623 503
1717 503
1717 525
4 12 27 0 0 8320 0 19 17 0 0 4
1605 497
1605 510
1708 510
1708 525
6 11 28 0 0 8320 0 19 17 0 0 4
1587 497
1587 517
1699 517
1699 525
8 10 29 0 0 8320 0 19 17 0 0 3
1569 497
1569 525
1690 525
0 1 3 0 0 0 0 0 17 54 0 3
1553 653
1663 653
1663 589
0 2 4 0 0 0 0 0 17 55 0 3
1573 644
1672 644
1672 589
0 3 5 0 0 0 0 0 17 56 0 3
1590 633
1681 633
1681 589
0 4 6 0 0 0 0 0 17 57 0 3
1609 626
1690 626
1690 589
1 0 2 0 0 0 0 23 0 0 47 3
1266 337
1266 359
1257 359
2 0 2 0 0 4224 0 23 0 0 48 2
1257 337
1257 373
3 1 2 0 0 0 0 23 18 0 0 3
1248 337
1248 373
1262 373
14 1 30 0 0 8320 0 19 22 0 0 4
1560 433
1560 390
1614 390
1614 341
13 2 31 0 0 12416 0 19 22 0 0 4
1578 433
1578 401
1605 401
1605 341
3 12 32 0 0 4224 0 22 19 0 0 2
1596 341
1596 433
4 11 33 0 0 4224 0 22 19 0 0 4
1587 341
1587 408
1614 408
1614 433
1 4 25 0 0 0 0 19 13 0 0 5
1632 497
1632 545
1461 545
1461 508
1394 508
10 9 3 0 0 128 0 8 19 0 0 8
1443 897
1443 909
1551 909
1551 690
1423 690
1423 653
1560 653
1560 497
11 7 4 0 0 128 0 8 19 0 0 8
1434 897
1434 918
1541 918
1541 694
1414 694
1414 644
1578 644
1578 497
12 5 5 0 0 128 0 8 19 0 0 10
1425 897
1425 937
1534 937
1534 704
1405 704
1405 666
1408 666
1408 633
1596 633
1596 497
13 3 6 0 0 128 0 8 19 0 0 8
1416 897
1416 949
1526 949
1526 710
1396 710
1396 626
1614 626
1614 497
1 2 34 0 0 4224 0 20 26 0 0 2
1600 68
1600 91
9 1 35 0 0 4224 0 21 26 0 0 2
1600 133
1600 127
13 1 36 0 0 12416 0 22 21 0 0 5
1560 271
1560 240
1580 240
1580 205
1579 205
12 2 37 0 0 12416 0 22 21 0 0 5
1569 271
1569 248
1586 248
1586 205
1585 205
11 3 38 0 0 12416 0 22 21 0 0 5
1578 271
1578 258
1592 258
1592 205
1591 205
4 10 39 0 0 16512 0 21 22 0 0 7
1597 205
1598 205
1598 209
1596 209
1596 264
1587 264
1587 271
5 9 40 0 0 16512 0 21 22 0 0 6
1603 205
1604 205
1604 212
1600 212
1600 271
1596 271
8 6 41 0 0 4224 0 22 21 0 0 5
1605 271
1605 216
1610 216
1610 205
1609 205
7 7 42 0 0 12416 0 21 22 0 0 4
1615 205
1615 203
1614 203
1614 271
1 2 43 0 0 4224 0 25 27 0 0 2
1252 64
1252 87
9 1 44 0 0 4224 0 24 27 0 0 2
1252 129
1252 123
13 1 45 0 0 12416 0 23 24 0 0 5
1212 267
1212 236
1232 236
1232 201
1231 201
12 2 46 0 0 12416 0 23 24 0 0 5
1221 267
1221 244
1238 244
1238 201
1237 201
11 3 47 0 0 12416 0 23 24 0 0 5
1230 267
1230 254
1244 254
1244 201
1243 201
4 10 48 0 0 16512 0 24 23 0 0 7
1249 201
1250 201
1250 205
1248 205
1248 260
1239 260
1239 267
5 9 49 0 0 16512 0 24 23 0 0 6
1255 201
1256 201
1256 208
1252 208
1252 267
1248 267
8 6 50 0 0 4224 0 23 24 0 0 5
1257 267
1257 212
1262 212
1262 201
1261 201
7 7 51 0 0 12416 0 24 23 0 0 4
1267 201
1267 199
1266 199
1266 267
3
-19 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 12
967 93 1091 122
975 100 1091 121
12 ASCII Keypad
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1877 125 1909 146
1884 132 1908 147
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1767 124 1799 145
1774 131 1798 146
3 MSB
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
