CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 50 3 80 9
0 71 1536 864
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 864
177209362 0
0
6 Title:
5 Name:
0
0
0
35
13 Logic Switch~
5 69 622 0 10 11
0 74 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 166 649 0 1 11
0 73
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 908 724 0 1 11
0 65
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 936 739 0 10 11
0 64 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V6
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 965 756 0 10 11
0 63 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V7
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 995 774 0 1 11
0 62
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V8
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 779 543 0 1 11
0 36
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V9
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 278 358 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 337 671 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3549 0 0
0
0
6 74LS47
187 780 287 0 14 29
0 4 3 5 6 75 76 15 14 13
12 11 10 9 77
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
3 U10
57 0 78 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
9 CA 7-Seg~
184 798 188 0 18 19
10 9 10 11 12 13 14 15 78 7
2 0 0 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9325 0 0
0
0
2 +V
167 798 103 0 1 3
0 8
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V14
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
2 +V
167 536 107 0 1 3
0 17
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V13
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3834 0 0
0
0
9 CA 7-Seg~
184 536 192 0 18 19
10 18 19 20 21 22 23 24 79 16
0 0 2 0 0 2 0 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3363 0 0
0
0
6 74LS47
187 518 291 0 14 29
0 32 31 30 28 80 81 24 23 22
21 20 19 18 82
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U4
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
7 Pulser~
4 32 565 0 10 12
0 83 84 85 35 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4718 0 0
0
0
9 2-In AND~
219 129 582 0 3 22
0 35 74 72
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3874 0 0
0
0
8 2-In OR~
219 208 597 0 3 22
0 72 73 34
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 3 0
1 U
6671 0 0
0
0
7 74LS273
150 655 703 0 18 37
0 61 27 45 46 47 48 49 50 51
52 71 70 69 68 4 3 5 6
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
2 U9
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
3789 0 0
0
0
7 Ground~
168 885 812 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4871 0 0
0
0
6 74LS83
105 815 828 0 14 29
0 4 3 5 6 65 64 63 62 2
57 58 59 60 67
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U8
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3750 0 0
0
0
6 74LS83
105 670 828 0 14 29
0 71 70 69 68 66 66 66 66 67
56 55 54 53 33
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U5
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
8778 0 0
0
0
2 +V
167 702 773 0 1 3
0 66
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
538 0 0
0
0
7 74LS157
122 683 565 0 14 29
0 36 44 60 43 59 42 58 41 57
2 52 51 50 49
0
0 0 13040 270
7 74LS157
-24 -60 25 -52
2 U1
54 0 68 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
6843 0 0
0
0
7 74LS157
122 555 562 0 14 29
0 36 40 53 39 54 38 55 37 56
2 48 47 46 45
0
0 0 13040 270
7 74LS157
-24 -60 25 -52
2 U2
54 0 68 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3136 0 0
0
0
10 Ascii Key~
169 678 451 0 11 12
0 44 43 42 41 86 87 88 89 0
0 53
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
5950 0 0
0
0
10 Ascii Key~
169 544 452 0 11 12
0 40 39 38 37 90 91 92 93 0
0 49
0
0 0 4656 0
0
4 KBD2
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
5670 0 0
0
0
9 2-In AND~
219 288 645 0 3 22
0 34 33 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
6828 0 0
0
0
6 74LS93
109 360 377 0 8 17
0 29 29 25 28 32 31 30 28
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
2 U3
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
6735 0 0
0
0
7 Ground~
168 493 529 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8365 0 0
0
0
7 Ground~
168 623 541 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4132 0 0
0
0
8 2-In OR~
219 375 661 0 3 22
0 25 26 27
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
4551 0 0
0
0
2 +V
167 584 674 0 1 3
0 61
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V12
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3635 0 0
0
0
9 Resistor~
219 799 127 0 4 5
0 7 8 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3973 0 0
0
0
9 Resistor~
219 537 131 0 4 5
0 16 17 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3851 0 0
0
0
88
2 0 3 0 0 4224 0 10 0 0 79 4
812 324
812 691
778 691
778 751
0 1 4 0 0 12416 0 0 10 78 0 4
771 757
771 684
821 684
821 324
0 3 5 0 0 12416 0 0 10 80 0 4
786 745
786 695
803 695
803 324
4 0 6 0 0 4224 0 10 0 0 81 2
794 324
794 740
1 9 7 0 0 8336 0 34 11 0 0 3
799 145
798 145
798 152
1 2 8 0 0 4240 0 12 34 0 0 3
798 112
798 109
799 109
1 13 9 0 0 4240 0 11 10 0 0 4
777 224
777 244
767 244
767 254
2 12 10 0 0 4240 0 11 10 0 0 4
783 224
783 249
776 249
776 254
3 11 11 0 0 4240 0 11 10 0 0 3
789 224
789 254
785 254
4 10 12 0 0 8336 0 11 10 0 0 3
795 224
794 224
794 254
5 9 13 0 0 8336 0 11 10 0 0 3
801 224
803 224
803 254
6 8 14 0 0 12432 0 11 10 0 0 4
807 224
807 237
812 237
812 254
7 7 15 0 0 12432 0 11 10 0 0 4
813 224
813 234
821 234
821 254
1 9 16 0 0 8320 0 35 14 0 0 3
537 149
536 149
536 156
1 2 17 0 0 4224 0 13 35 0 0 3
536 116
536 113
537 113
1 13 18 0 0 4224 0 14 15 0 0 4
515 228
515 248
505 248
505 258
2 12 19 0 0 4224 0 14 15 0 0 4
521 228
521 253
514 253
514 258
3 11 20 0 0 4224 0 14 15 0 0 3
527 228
527 258
523 258
4 10 21 0 0 8320 0 14 15 0 0 3
533 228
532 228
532 258
5 9 22 0 0 8320 0 14 15 0 0 3
539 228
541 228
541 258
6 8 23 0 0 12416 0 14 15 0 0 4
545 228
545 241
550 241
550 258
7 7 24 0 0 12416 0 14 15 0 0 4
551 228
551 238
559 238
559 258
3 0 25 0 0 8320 0 29 0 0 27 3
322 386
316 386
316 645
1 0 26 0 0 4096 0 9 0 0 25 2
349 671
349 670
2 0 26 0 0 4224 0 32 0 0 0 2
362 670
345 670
3 2 27 0 0 4224 0 32 19 0 0 3
408 661
623 661
623 676
3 1 25 0 0 0 0 28 32 0 0 4
309 645
353 645
353 652
362 652
4 0 28 0 0 8192 0 29 0 0 30 4
322 395
322 411
402 411
402 395
1 0 29 0 0 4096 0 8 0 0 34 2
290 358
290 357
8 4 28 0 0 4224 0 29 15 0 0 3
392 395
532 395
532 328
7 3 30 0 0 4224 0 29 15 0 0 3
392 386
541 386
541 328
6 2 31 0 0 4224 0 29 15 0 0 3
392 377
550 377
550 328
5 1 32 0 0 4224 0 29 15 0 0 3
392 368
559 368
559 328
0 1 29 0 0 4224 0 0 29 0 0 3
286 357
328 357
328 368
1 2 29 0 0 0 0 29 29 0 0 2
328 368
328 377
1 10 2 0 0 4096 0 30 25 0 0 3
493 523
509 523
509 529
1 10 2 0 0 0 0 31 24 0 0 4
623 535
623 527
637 527
637 532
2 14 33 0 0 8320 0 28 22 0 0 4
264 654
264 908
713 908
713 862
3 1 34 0 0 8320 0 18 28 0 0 3
241 597
264 597
264 636
4 1 35 0 0 4224 0 16 17 0 0 3
62 565
105 565
105 573
0 1 36 0 0 4096 0 0 7 66 0 3
717 523
767 523
767 543
8 4 37 0 0 4224 0 25 27 0 0 4
527 535
527 489
547 489
547 476
3 6 38 0 0 12416 0 27 25 0 0 4
553 476
553 494
545 494
545 535
2 4 39 0 0 4224 0 27 25 0 0 4
559 476
559 531
563 531
563 535
1 2 40 0 0 8320 0 27 25 0 0 3
565 476
581 476
581 535
4 8 41 0 0 12416 0 26 24 0 0 4
681 475
681 488
655 488
655 538
3 6 42 0 0 12416 0 26 24 0 0 4
687 475
687 494
673 494
673 538
2 4 43 0 0 8320 0 26 24 0 0 3
693 475
691 475
691 538
1 2 44 0 0 8320 0 26 24 0 0 3
699 475
709 475
709 538
14 3 45 0 0 8320 0 25 19 0 0 4
518 599
518 656
632 656
632 676
13 4 46 0 0 8320 0 25 19 0 0 4
536 599
536 650
641 650
641 676
12 5 47 0 0 8320 0 25 19 0 0 4
554 599
554 646
650 646
650 676
11 6 48 0 0 8320 0 25 19 0 0 4
572 599
572 643
659 643
659 676
14 7 49 0 0 12416 0 24 19 0 0 4
646 602
646 638
668 638
668 676
13 8 50 0 0 12416 0 24 19 0 0 4
664 602
664 633
677 633
677 676
12 9 51 0 0 4224 0 24 19 0 0 3
682 602
682 676
686 676
11 10 52 0 0 4224 0 24 19 0 0 3
700 602
700 676
695 676
13 3 53 0 0 12416 0 22 25 0 0 6
686 862
686 898
453 898
453 500
572 500
572 535
12 5 54 0 0 12416 0 22 25 0 0 6
677 862
677 891
460 891
460 504
554 504
554 535
7 11 55 0 0 12416 0 25 22 0 0 6
536 535
536 508
468 508
468 885
668 885
668 862
9 10 56 0 0 12416 0 25 22 0 0 6
518 535
518 511
481 511
481 869
659 869
659 862
10 9 57 0 0 12416 0 21 24 0 0 6
804 862
804 898
1043 898
1043 500
646 500
646 538
11 7 58 0 0 12416 0 21 24 0 0 6
813 862
813 890
1028 890
1028 504
664 504
664 538
12 5 59 0 0 12416 0 21 24 0 0 6
822 862
822 884
1023 884
1023 507
682 507
682 538
13 3 60 0 0 12416 0 21 24 0 0 6
831 862
831 877
1015 877
1015 518
700 518
700 538
1 1 36 0 0 8320 0 25 24 0 0 4
590 535
590 523
718 523
718 538
1 1 61 0 0 4224 0 19 33 0 0 4
614 670
583 670
583 683
584 683
8 1 62 0 0 8320 0 21 6 0 0 3
840 798
840 774
983 774
7 1 63 0 0 8320 0 21 5 0 0 3
831 798
831 756
953 756
6 1 64 0 0 8320 0 21 4 0 0 3
822 798
822 739
924 739
5 1 65 0 0 8320 0 21 3 0 0 3
813 798
813 724
896 724
0 1 66 0 0 4224 0 0 23 73 0 4
689 798
689 780
702 780
702 782
7 8 66 0 0 0 0 22 22 0 0 2
686 798
695 798
6 7 66 0 0 0 0 22 22 0 0 2
677 798
686 798
5 6 66 0 0 0 0 22 22 0 0 2
668 798
677 798
9 1 2 0 0 4224 0 21 20 0 0 3
858 798
885 798
885 806
9 14 67 0 0 12416 0 22 21 0 0 5
713 798
747 798
747 869
858 869
858 862
15 1 4 0 0 0 0 19 21 0 0 4
668 740
668 757
777 757
777 798
16 2 3 0 0 128 0 19 21 0 0 4
677 740
677 751
786 751
786 798
17 3 5 0 0 0 0 19 21 0 0 4
686 740
686 745
795 745
795 798
18 4 6 0 0 0 0 19 21 0 0 3
695 740
804 740
804 798
14 4 68 0 0 4224 0 19 22 0 0 2
659 740
659 798
13 3 69 0 0 4224 0 19 22 0 0 2
650 740
650 798
12 2 70 0 0 4224 0 19 22 0 0 2
641 740
641 798
11 1 71 0 0 4224 0 19 22 0 0 2
632 740
632 798
3 1 72 0 0 4224 0 17 18 0 0 4
150 582
185 582
185 588
195 588
2 1 73 0 0 8320 0 18 2 0 0 4
195 606
185 606
185 649
178 649
2 1 74 0 0 8320 0 17 1 0 0 4
105 591
92 591
92 622
81 622
4
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
269 686 402 723
282 696 402 721
10 select clk
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
827 529 996 566
841 539 997 564
13 select contro
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
49 515 218 552
62 525 218 550
13 Clock control
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
107 655 264 692
116 662 260 687
12 Manual clock
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
