CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
500 110 1 80 9
0 76 1536 869
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 76 1536 869
143654930 0
0
6 Title:
5 Name:
0
0
0
32
13 Logic Switch~
5 1705 843 0 1 11
0 33
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 1639 809 0 1 11
0 36
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 1557 781 0 1 11
0 35
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V9
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 1504 755 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V8
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
9 Inverter~
13 1086 752 0 2 22
0 3 4
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U10E
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 6 0
1 U
5394 0 0
0
0
9 2-In AND~
219 1441 562 0 3 22
0 6 7 5
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U8A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1979603804
65 0 0 0 4 1 9 0
1 U
7734 0 0
0
0
8 2-In OR~
219 1398 604 0 3 22
0 9 8 6
0
0 0 624 90
6 74LS32
-21 -24 21 -16
3 U6B
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 8 0
1 U
9914 0 0
0
0
8 2-In OR~
219 1390 535 0 3 22
0 10 5 22
0
0 0 624 90
6 74LS32
-21 -24 21 -16
3 U6A
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1459510143
65 0 0 0 4 1 8 0
1 U
3747 0 0
0
0
7 Buffer~
58 877 719 0 2 22
0 13 12
0
0 0 624 270
4 4050
-14 -19 14 -11
4 U11D
14 -5 42 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 4 7 0
1 U
3549 0 0
0
0
7 Buffer~
58 876 797 0 2 22
0 11 14
0
0 0 624 270
4 4050
-14 -19 14 -11
4 U11C
14 -5 42 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 3 7 0
1 U
7931 0 0
0
0
7 Buffer~
58 877 755 0 2 22
0 12 11
0
0 0 624 270
4 4050
-14 -19 14 -11
4 U11B
14 -5 42 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 2 7 0
1 U
9325 0 0
0
0
9 Inverter~
13 1105 733 0 2 22
0 17 21
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U10D
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 6 0
1 U
8903 0 0
0
0
7 Buffer~
58 1081 277 0 2 22
0 15 16
0
0 0 624 0
4 4050
-14 -19 14 -11
4 U11A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 7 0
1 U
3834 0 0
0
0
9 Inverter~
13 1123 714 0 2 22
0 18 20
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U10C
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 6 0
1 U
3363 0 0
0
0
9 4-In AND~
219 1045 738 0 5 22
0 19 20 21 4 13
0
0 0 624 512
6 74LS21
-21 -28 21 -20
3 U5A
-13 -28 8 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 2130598743
65 0 0 0 2 1 5 0
1 U
7668 0 0
0
0
7 Pulser~
4 991 858 0 10 12
0 54 55 15 56 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4718 0 0
0
0
6 74LS93
109 1078 832 0 8 17
0 14 57 15 3 19 18 17 3
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
2 U4
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
7 Ground~
168 1331 738 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6671 0 0
0
0
7 Ground~
168 1543 526 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3789 0 0
0
0
7 Ground~
168 1817 659 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4871 0 0
0
0
6 74LS83
105 1803 552 0 14 29
0 7 8 9 27 2 28 28 2 2
26 25 24 23 58
0
0 0 13040 90
7 74LS83A
-24 -60 25 -52
2 U9
57 -3 71 5
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3750 0 0
0
0
7 Ground~
168 1262 379 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8778 0 0
0
0
7 74LS157
122 1593 462 0 14 29
0 22 23 27 24 9 25 8 26 7
2 32 31 30 29
0
0 0 13040 602
7 74LS157
-24 -60 25 -52
2 U7
54 -6 68 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
538 0 0
0
0
6 74LS83
105 1412 696 0 14 29
0 34 35 36 33 19 18 17 3 2
7 8 9 27 10
0
0 0 13040 602
7 74LS83A
-24 -60 25 -52
2 U3
57 -3 71 5
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6843 0 0
0
0
2 +V
167 1600 59 0 1 3
0 28
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3136 0 0
0
0
9 CA 7-Seg~
184 1600 169 0 18 19
10 38 39 40 41 42 43 44 59 37
2 2 2 0 0 2 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5950 0 0
0
0
6 74LS47
187 1573 304 0 14 29
0 29 30 31 32 60 61 44 43 42
41 40 39 38 16
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
6 74LS47
187 1225 300 0 14 29
0 2 2 2 22 62 63 53 52 51
50 49 48 47 16
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U2
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6828 0 0
0
0
9 CA 7-Seg~
184 1252 165 0 18 19
10 47 48 49 50 51 52 53 64 46
2 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6735 0 0
0
0
2 +V
167 1252 55 0 1 3
0 45
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8365 0 0
0
0
9 Resistor~
219 1600 109 0 4 5
0 37 28 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 1252 105 0 4 5
0 46 45 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
78
1 0 3 0 0 8192 0 5 0 0 56 3
1107 752
1117 752
1117 850
4 2 4 0 0 4224 0 15 5 0 0 2
1065 752
1071 752
2 3 5 0 0 16512 0 8 6 0 0 5
1402 551
1402 556
1411 556
1411 538
1440 538
3 1 6 0 0 4224 0 7 6 0 0 5
1401 574
1421 574
1421 586
1431 586
1431 583
0 2 7 0 0 4096 0 0 6 48 0 3
1452 653
1452 583
1449 583
2 0 8 0 0 8192 0 7 0 0 49 3
1410 620
1420 620
1420 644
1 0 9 0 0 4096 0 7 0 0 50 3
1392 620
1392 642
1408 642
14 1 10 0 0 4224 0 24 8 0 0 4
1369 666
1369 554
1384 554
1384 551
2 1 11 0 0 8320 0 11 10 0 0 3
877 770
876 770
876 782
2 1 12 0 0 4224 0 9 11 0 0 2
877 734
877 740
1 5 13 0 0 4224 0 9 15 0 0 4
877 704
995 704
995 738
1020 738
2 1 14 0 0 4224 0 10 17 0 0 4
876 812
1036 812
1036 823
1046 823
0 1 15 0 0 4224 0 0 13 21 0 3
1015 842
1015 277
1066 277
0 14 16 0 0 8320 0 0 27 15 0 6
1145 277
1145 393
1488 393
1488 264
1533 264
1533 277
2 14 16 0 0 0 0 13 28 0 0 4
1096 277
1145 277
1145 273
1185 273
1 0 17 0 0 4096 0 12 0 0 55 2
1126 733
1126 841
1 0 18 0 0 4096 0 14 0 0 54 2
1144 714
1144 832
1 0 19 0 0 12288 0 15 0 0 53 4
1065 725
1065 690
1196 690
1196 823
2 2 20 0 0 12416 0 15 14 0 0 4
1065 734
1070 734
1070 714
1108 714
3 2 21 0 0 12416 0 15 12 0 0 4
1065 743
1075 743
1075 733
1090 733
3 3 15 0 0 128 0 16 17 0 0 3
1015 849
1015 841
1040 841
0 4 3 0 0 0 0 0 17 56 0 4
1123 850
1123 892
1040 892
1040 850
1 0 2 0 0 4096 0 18 0 0 24 2
1331 732
1331 730
9 0 2 0 0 4096 0 24 0 0 0 3
1369 730
1331 730
1331 736
10 1 2 0 0 0 0 23 19 0 0 4
1547 499
1547 514
1543 514
1543 520
4 0 22 0 0 8320 0 28 0 0 47 4
1239 337
1239 459
1417 459
1417 508
2 13 23 0 0 8320 0 23 21 0 0 4
1619 493
1619 503
1819 503
1819 522
4 12 24 0 0 8320 0 23 21 0 0 4
1601 493
1601 510
1810 510
1810 522
6 11 25 0 0 8320 0 23 21 0 0 4
1583 493
1583 517
1801 517
1801 522
8 10 26 0 0 8320 0 23 21 0 0 3
1565 493
1565 522
1792 522
0 1 7 0 0 4224 0 0 21 48 0 3
1553 653
1765 653
1765 586
0 2 8 0 0 4224 0 0 21 49 0 3
1573 644
1774 644
1774 586
0 3 9 0 0 4224 0 0 21 50 0 3
1590 633
1783 633
1783 586
0 4 27 0 0 4096 0 0 21 51 0 3
1609 626
1792 626
1792 586
6 0 28 0 0 4096 0 21 0 0 36 3
1810 586
1810 604
1819 604
0 7 28 0 0 8320 0 0 21 61 0 5
1600 82
2007 82
2007 604
1819 604
1819 586
9 0 2 0 0 0 0 21 0 0 38 3
1846 586
1846 624
1828 624
8 1 2 0 0 4224 0 21 20 0 0 3
1828 586
1828 653
1817 653
5 1 2 0 0 0 0 21 20 0 0 3
1801 586
1801 653
1817 653
1 0 2 0 0 0 0 28 0 0 41 3
1266 337
1266 359
1257 359
2 0 2 0 0 0 0 28 0 0 42 2
1257 337
1257 373
3 1 2 0 0 0 0 28 22 0 0 3
1248 337
1248 373
1262 373
14 1 29 0 0 8320 0 23 27 0 0 4
1556 429
1556 390
1614 390
1614 341
13 2 30 0 0 12416 0 23 27 0 0 4
1574 429
1574 401
1605 401
1605 341
3 12 31 0 0 4224 0 27 23 0 0 4
1596 341
1596 422
1592 422
1592 429
4 11 32 0 0 4224 0 27 23 0 0 4
1587 341
1587 408
1610 408
1610 429
1 3 22 0 0 0 0 23 8 0 0 6
1628 493
1628 545
1461 545
1461 508
1393 508
1393 505
10 9 7 0 0 0 0 24 23 0 0 4
1423 666
1423 653
1556 653
1556 493
11 7 8 0 0 0 0 24 23 0 0 4
1414 666
1414 644
1574 644
1574 493
12 5 9 0 0 0 0 24 23 0 0 5
1405 666
1408 666
1408 633
1592 633
1592 493
13 3 27 0 0 8320 0 24 23 0 0 4
1396 666
1396 626
1610 626
1610 493
1 0 33 0 0 0 0 1 0 0 60 2
1693 843
1693 843
5 5 19 0 0 12416 0 17 24 0 0 5
1110 823
1206 823
1206 762
1414 762
1414 730
6 6 18 0 0 12416 0 17 24 0 0 5
1110 832
1223 832
1223 813
1405 813
1405 730
7 7 17 0 0 12416 0 17 24 0 0 5
1110 841
1181 841
1181 865
1396 865
1396 730
8 8 3 0 0 12416 0 17 24 0 0 5
1110 850
1160 850
1160 915
1387 915
1387 730
1 1 34 0 0 8320 0 24 4 0 0 4
1450 730
1450 756
1492 756
1492 755
2 1 35 0 0 8320 0 24 3 0 0 3
1441 730
1441 781
1545 781
3 1 36 0 0 8320 0 24 2 0 0 4
1432 730
1432 808
1627 808
1627 809
4 0 33 0 0 8320 0 24 0 0 0 3
1423 730
1423 843
1699 843
1 2 28 0 0 0 0 25 31 0 0 2
1600 68
1600 91
9 1 37 0 0 4224 0 26 31 0 0 2
1600 133
1600 127
13 1 38 0 0 12416 0 27 26 0 0 5
1560 271
1560 240
1580 240
1580 205
1579 205
12 2 39 0 0 12416 0 27 26 0 0 5
1569 271
1569 248
1586 248
1586 205
1585 205
11 3 40 0 0 12416 0 27 26 0 0 5
1578 271
1578 258
1592 258
1592 205
1591 205
4 10 41 0 0 16512 0 26 27 0 0 7
1597 205
1598 205
1598 209
1596 209
1596 264
1587 264
1587 271
5 9 42 0 0 16512 0 26 27 0 0 6
1603 205
1604 205
1604 212
1600 212
1600 271
1596 271
8 6 43 0 0 4224 0 27 26 0 0 5
1605 271
1605 216
1610 216
1610 205
1609 205
7 7 44 0 0 12416 0 26 27 0 0 4
1615 205
1615 203
1614 203
1614 271
1 2 45 0 0 4224 0 30 32 0 0 2
1252 64
1252 87
9 1 46 0 0 4224 0 29 32 0 0 2
1252 129
1252 123
13 1 47 0 0 12416 0 28 29 0 0 5
1212 267
1212 236
1232 236
1232 201
1231 201
12 2 48 0 0 12416 0 28 29 0 0 5
1221 267
1221 244
1238 244
1238 201
1237 201
11 3 49 0 0 12416 0 28 29 0 0 5
1230 267
1230 254
1244 254
1244 201
1243 201
4 10 50 0 0 16512 0 29 28 0 0 7
1249 201
1250 201
1250 205
1248 205
1248 260
1239 260
1239 267
5 9 51 0 0 16512 0 29 28 0 0 6
1255 201
1256 201
1256 208
1252 208
1252 267
1248 267
8 6 52 0 0 4224 0 28 29 0 0 5
1257 267
1257 212
1262 212
1262 201
1261 201
7 7 53 0 0 12416 0 29 28 0 0 4
1267 201
1267 199
1266 199
1266 267
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
