CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1020 230 2 200 9
0 76 1534 869
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 76 1534 869
143654930 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 1263 277 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
6 74LS83
105 1554 430 0 14 29
0 16 15 14 13 5 6 7 8 2
21 20 19 18 22
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
3 U11
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
4441 0 0
0
0
14 Logic Display~
6 1559 511 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 1586 511 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 1532 512 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 1506 512 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 1478 514 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
7 Buffer~
58 1102 355 0 2 22
0 4 3
0
0 0 624 270
4 4050
-14 -19 14 -11
4 U12A
14 -5 42 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 5 0
1 U
3747 0 0
0
0
7 74LS273
150 1329 317 0 18 37
0 17 3 5 6 7 8 9 10 11
12 16 15 14 13 5 6 7 8
0
0 0 13040 0
7 74LS273
-24 -60 25 -52
3 U10
-11 -61 10 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
10 Ascii Key~
169 1144 285 0 11 12
0 12 11 10 9 23 24 25 4 0
0 56
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
7931 0 0
0
0
7 Ground~
168 1479 407 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
25
2 2 3 0 0 8320 0 8 9 0 0 5
1102 370
1102 404
1246 404
1246 290
1297 290
8 1 4 0 0 4224 0 10 8 0 0 4
1123 309
1123 335
1102 335
1102 340
0 3 5 0 0 8192 0 0 9 15 0 5
1405 335
1405 413
1260 413
1260 299
1297 299
0 4 6 0 0 8192 0 0 9 14 0 5
1396 344
1396 400
1271 400
1271 308
1297 308
0 5 7 0 0 8192 0 0 9 13 0 5
1384 353
1384 388
1278 388
1278 317
1297 317
0 6 8 0 0 8192 0 0 9 12 0 5
1373 362
1373 379
1289 379
1289 326
1297 326
4 7 9 0 0 8320 0 10 9 0 0 3
1147 309
1147 335
1297 335
3 8 10 0 0 8320 0 10 9 0 0 3
1153 309
1153 344
1297 344
2 9 11 0 0 8320 0 10 9 0 0 3
1159 309
1159 353
1297 353
1 10 12 0 0 8320 0 10 9 0 0 3
1165 309
1165 362
1297 362
9 1 2 0 0 8320 0 2 11 0 0 4
1511 400
1511 372
1479 372
1479 401
18 8 8 0 0 4224 0 9 2 0 0 3
1361 362
1529 362
1529 400
17 7 7 0 0 4224 0 9 2 0 0 3
1361 353
1538 353
1538 400
16 6 6 0 0 4224 0 9 2 0 0 3
1361 344
1547 344
1547 400
15 5 5 0 0 4224 0 9 2 0 0 3
1361 335
1556 335
1556 400
14 4 13 0 0 4224 0 9 2 0 0 3
1361 326
1565 326
1565 400
13 3 14 0 0 4224 0 9 2 0 0 3
1361 317
1574 317
1574 400
12 2 15 0 0 4224 0 9 2 0 0 3
1361 308
1583 308
1583 400
11 1 16 0 0 4224 0 9 2 0 0 3
1361 299
1592 299
1592 400
1 1 17 0 0 4224 0 1 9 0 0 3
1275 277
1291 277
1291 281
13 1 18 0 0 8320 0 2 4 0 0 6
1538 464
1538 485
1606 485
1606 535
1586 535
1586 529
12 1 19 0 0 8320 0 2 3 0 0 6
1547 464
1547 479
1631 479
1631 541
1559 541
1559 529
11 1 20 0 0 16512 0 2 5 0 0 6
1556 464
1556 473
1646 473
1646 555
1532 555
1532 530
10 1 21 0 0 12416 0 2 6 0 0 5
1565 464
1659 464
1659 568
1506 568
1506 530
14 1 22 0 0 12416 0 2 7 0 0 6
1511 464
1511 472
1464 472
1464 537
1478 537
1478 532
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
