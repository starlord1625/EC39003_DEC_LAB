CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1120 20 5 120 9
0 71 1536 864
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 864
143654930 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 1449 270 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 1474 312 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 1789 426 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 1326 584 0 1 11
0 45
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 1183 557 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 1369 453 0 1 11
0 46
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
9 CC 7-Seg~
183 2320 116 0 18 19
10 12 13 14 15 16 17 18 54 4
0 1 1 0 0 0 0 2 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP9
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
9914 0 0
0
0
9 CC 7-Seg~
183 2261 115 0 18 19
10 12 13 14 15 16 17 18 55 5
0 1 1 0 0 0 0 2 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP8
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3747 0 0
0
0
9 CC 7-Seg~
183 2198 114 0 18 19
10 12 13 14 15 16 17 18 56 6
0 1 1 0 0 0 0 2 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP7
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3549 0 0
0
0
9 CC 7-Seg~
183 2134 112 0 17 19
10 12 13 14 15 16 17 18 57 7
0 1 1 0 0 0 0 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
7931 0 0
0
0
9 CC 7-Seg~
183 2072 112 0 18 19
10 12 13 14 15 16 17 18 58 8
0 1 1 0 0 0 0 2 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP5
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
9325 0 0
0
0
9 CC 7-Seg~
183 2007 111 0 18 19
10 12 13 14 15 16 17 18 59 9
0 1 1 0 0 0 0 2 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
8903 0 0
0
0
9 CC 7-Seg~
183 1939 112 0 18 19
10 12 13 14 15 16 17 18 60 10
0 1 1 0 0 0 0 2 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3834 0 0
0
0
6 74LS48
188 1735 343 0 14 29
0 22 21 20 19 61 3 18 17 16
15 14 13 12 3
0
0 0 13040 0
6 74LS48
-21 -60 21 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3363 0 0
0
0
7 74LS138
19 1549 335 0 14 29
0 25 26 27 24 23 23 4 5 6
7 8 9 10 11
0
0 0 13296 692
7 74LS138
-25 -62 24 -54
2 U8
-7 -72 7 -64
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
9 CC 7-Seg~
183 1857 112 0 18 19
10 12 13 14 15 16 17 18 65 11
0 1 1 0 0 0 0 2 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
4718 0 0
0
0
7 Ground~
168 1521 442 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3874 0 0
0
0
7 Ground~
168 1652 431 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
7 Ground~
168 1922 462 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3789 0 0
0
0
8 2-In OR~
219 1368 532 0 3 22
0 44 45 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1330618039
65 0 0 0 4 1 3 0
1 U
4871 0 0
0
0
7 Pulser~
4 1200 502 0 10 12
0 66 67 42 68 0 0 5 5 3
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3750 0 0
0
0
9 2-In AND~
219 1280 530 0 3 22
0 42 43 44
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
8778 0 0
0
0
6 74LS93
109 1457 507 0 8 17
0 46 46 69 3 25 26 27 70
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
2 U5
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
538 0 0
0
0
7 Buffer~
58 1980 464 0 2 22
0 53 52
0
0 0 624 180
4 4050
-14 -19 14 -11
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
6843 0 0
0
0
10 Ascii Key~
169 2075 431 0 11 12
0 48 49 50 51 71 72 73 53 0
0 49
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3136 0 0
0
0
7 74LS173
129 1843 481 0 14 29
0 2 2 2 52 51 50 49 48 47
47 22 21 20 19
0
0 0 13040 512
7 74LS173
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
5950 0 0
0
0
6 1K RAM
79 1589 472 0 20 41
0 2 2 2 2 2 2 2 25 26
27 74 75 76 77 22 21 20 19 2
47
0
0 0 13040 0
5 RAM1K
-17 -19 18 -11
2 U1
-7 -70 7 -62
0
15 DVCC=22;DGND=11
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
119
0 0 3 0 0 8320 0 0 0 2 90 4
1738 415
1738 570
1413 570
1413 532
6 14 3 0 0 0 0 14 14 0 0 4
1703 388
1703 415
1767 415
1767 388
7 9 4 0 0 12416 0 15 7 0 0 5
1587 354
1634 354
1634 65
2320 65
2320 74
8 9 5 0 0 12416 0 15 8 0 0 5
1587 345
1628 345
1628 53
2261 53
2261 73
9 9 6 0 0 12416 0 15 9 0 0 5
1587 336
1623 336
1623 44
2198 44
2198 72
10 9 7 0 0 12416 0 15 10 0 0 5
1587 327
1619 327
1619 38
2134 38
2134 70
11 9 8 0 0 12416 0 15 11 0 0 5
1587 318
1613 318
1613 33
2072 33
2072 70
12 9 9 0 0 12416 0 15 12 0 0 5
1587 309
1608 309
1608 25
2007 25
2007 69
13 9 10 0 0 12416 0 15 13 0 0 5
1587 300
1601 300
1601 20
1939 20
1939 70
14 9 11 0 0 8320 0 15 16 0 0 5
1587 291
1596 291
1596 13
1857 13
1857 70
1 0 12 0 0 4112 0 7 0 0 68 2
2299 152
2299 223
2 0 13 0 0 4112 0 7 0 0 69 2
2305 152
2305 214
3 0 14 0 0 4112 0 7 0 0 70 2
2311 152
2311 204
4 0 15 0 0 4112 0 7 0 0 71 2
2317 152
2317 193
5 0 16 0 0 4112 0 7 0 0 67 2
2323 152
2323 185
6 0 17 0 0 4112 0 7 0 0 72 2
2329 152
2329 176
7 0 18 0 0 4112 0 7 0 0 73 2
2335 152
2335 167
1 0 12 0 0 4096 0 8 0 0 68 2
2240 151
2240 223
2 0 13 0 0 4096 0 8 0 0 69 2
2246 151
2246 214
3 0 14 0 0 4096 0 8 0 0 70 2
2252 151
2252 204
4 0 15 0 0 4096 0 8 0 0 71 2
2258 151
2258 193
5 0 16 0 0 4096 0 8 0 0 67 2
2264 151
2264 185
6 0 17 0 0 4096 0 8 0 0 72 2
2270 151
2270 176
7 0 18 0 0 4096 0 8 0 0 73 2
2276 151
2276 167
1 0 12 0 0 4096 0 9 0 0 68 2
2177 150
2177 223
2 0 13 0 0 4096 0 9 0 0 69 2
2183 150
2183 214
3 0 14 0 0 4096 0 9 0 0 70 2
2189 150
2189 204
4 0 15 0 0 4096 0 9 0 0 71 2
2195 150
2195 193
5 0 16 0 0 4096 0 9 0 0 67 2
2201 150
2201 185
6 0 17 0 0 4096 0 9 0 0 72 2
2207 150
2207 176
7 0 18 0 0 4096 0 9 0 0 73 2
2213 150
2213 167
1 0 12 0 0 4096 0 10 0 0 68 2
2113 148
2113 223
2 0 13 0 0 4096 0 10 0 0 69 2
2119 148
2119 214
3 0 14 0 0 4096 0 10 0 0 70 2
2125 148
2125 204
4 0 15 0 0 4096 0 10 0 0 71 2
2131 148
2131 193
5 0 16 0 0 4096 0 10 0 0 67 2
2137 148
2137 185
6 0 17 0 0 4096 0 10 0 0 72 2
2143 148
2143 176
7 0 18 0 0 4096 0 10 0 0 73 2
2149 148
2149 167
1 0 12 0 0 0 0 11 0 0 68 2
2051 148
2051 223
2 0 13 0 0 0 0 11 0 0 69 2
2057 148
2057 214
3 0 14 0 0 0 0 11 0 0 70 2
2063 148
2063 204
4 0 15 0 0 0 0 11 0 0 71 2
2069 148
2069 193
5 0 16 0 0 0 0 11 0 0 67 2
2075 148
2075 185
6 0 17 0 0 0 0 11 0 0 72 2
2081 148
2081 176
7 0 18 0 0 0 0 11 0 0 73 2
2087 148
2087 167
1 0 12 0 0 4096 0 12 0 0 68 2
1986 147
1986 223
2 0 13 0 0 4096 0 12 0 0 69 2
1992 147
1992 214
3 0 14 0 0 4096 0 12 0 0 70 2
1998 147
1998 204
4 0 15 0 0 4096 0 12 0 0 71 2
2004 147
2004 193
5 0 16 0 0 4096 0 12 0 0 67 2
2010 147
2010 185
6 0 17 0 0 4096 0 12 0 0 72 2
2016 147
2016 176
7 0 18 0 0 4096 0 12 0 0 73 2
2022 147
2022 167
1 0 12 0 0 0 0 13 0 0 68 2
1918 148
1918 223
2 0 13 0 0 0 0 13 0 0 69 2
1924 148
1924 214
3 0 14 0 0 0 0 13 0 0 70 2
1930 148
1930 204
4 0 15 0 0 0 0 13 0 0 71 2
1936 148
1936 193
5 0 16 0 0 0 0 13 0 0 67 2
1942 148
1942 185
6 0 17 0 0 0 0 13 0 0 72 2
1948 148
1948 176
7 0 18 0 0 0 0 13 0 0 73 2
1954 148
1954 167
1 0 12 0 0 0 0 16 0 0 68 2
1836 148
1836 223
2 0 13 0 0 0 0 16 0 0 69 2
1842 148
1842 214
3 0 14 0 0 0 0 16 0 0 70 2
1848 148
1848 204
4 0 15 0 0 0 0 16 0 0 71 2
1854 148
1854 193
5 0 16 0 0 0 0 16 0 0 67 2
1860 148
1860 185
6 0 17 0 0 0 0 16 0 0 72 2
1866 148
1866 176
7 0 18 0 0 0 0 16 0 0 73 2
1872 148
1872 167
9 0 16 0 0 12416 0 14 0 0 0 4
1767 325
1789 325
1789 185
2811 185
13 0 12 0 0 12416 0 14 0 0 0 4
1767 361
1825 361
1825 223
2802 223
12 0 13 0 0 12416 0 14 0 0 0 4
1767 352
1817 352
1817 214
2809 214
11 0 14 0 0 12416 0 14 0 0 0 4
1767 343
1806 343
1806 204
2812 204
10 0 15 0 0 12416 0 14 0 0 0 4
1767 334
1797 334
1797 193
2813 193
8 0 17 0 0 12416 0 14 0 0 0 4
1767 316
1784 316
1784 176
2813 176
7 0 18 0 0 12416 0 14 0 0 0 4
1767 307
1774 307
1774 167
2810 167
4 0 19 0 0 8192 0 14 0 0 105 3
1703 334
1684 334
1684 517
3 0 20 0 0 8192 0 14 0 0 106 3
1703 325
1675 325
1675 508
2 0 21 0 0 8192 0 14 0 0 107 3
1703 316
1670 316
1670 499
1 0 22 0 0 8192 0 14 0 0 108 3
1703 307
1664 307
1664 490
1 0 23 0 0 0 0 1 0 0 79 2
1461 270
1461 270
0 0 23 0 0 8320 0 0 0 81 0 3
1499 291
1499 270
1458 270
1 0 24 0 0 0 0 2 0 0 82 2
1486 312
1486 312
6 5 23 0 0 0 0 15 15 0 0 4
1511 291
1498 291
1498 300
1511 300
0 4 24 0 0 4224 0 0 15 0 0 3
1483 312
1517 312
1517 309
1 0 25 0 0 8320 0 15 0 0 95 3
1517 354
1509 354
1509 498
2 0 26 0 0 8320 0 15 0 0 94 3
1517 345
1503 345
1503 508
3 0 27 0 0 8320 0 15 0 0 93 3
1517 336
1497 336
1497 517
3 1 42 0 0 8320 0 21 22 0 0 4
1224 493
1238 493
1238 521
1256 521
1 2 43 0 0 4224 0 5 22 0 0 4
1195 557
1238 557
1238 539
1256 539
3 1 44 0 0 8320 0 22 20 0 0 3
1301 530
1301 523
1355 523
2 1 45 0 0 8320 0 20 4 0 0 4
1355 541
1345 541
1345 584
1338 584
3 4 3 0 0 128 0 20 23 0 0 3
1401 532
1419 532
1419 525
0 1 46 0 0 8192 0 0 23 92 0 3
1415 497
1415 498
1425 498
1 2 46 0 0 8320 0 6 23 0 0 4
1381 453
1415 453
1415 507
1425 507
7 10 27 0 0 128 0 23 27 0 0 3
1489 516
1489 517
1557 517
6 9 26 0 0 128 0 23 27 0 0 3
1489 507
1489 508
1557 508
8 5 25 0 0 128 0 27 23 0 0 3
1557 499
1557 498
1489 498
2 0 2 0 0 4096 0 27 0 0 101 2
1557 445
1532 445
3 0 2 0 0 0 0 27 0 0 101 2
1557 454
1532 454
4 0 2 0 0 0 0 27 0 0 101 2
1557 463
1532 463
5 0 2 0 0 0 0 27 0 0 101 2
1557 472
1532 472
6 0 2 0 0 0 0 27 0 0 101 2
1557 481
1532 481
0 7 2 0 0 4224 0 0 27 102 0 3
1532 436
1532 490
1557 490
1 1 2 0 0 0 0 17 27 0 0 2
1521 436
1557 436
19 1 2 0 0 0 0 27 18 0 0 4
1627 436
1627 420
1652 420
1652 425
20 0 47 0 0 4224 0 27 0 0 110 2
1627 445
1801 445
18 14 19 0 0 4224 0 27 26 0 0 2
1621 517
1811 517
13 17 20 0 0 4224 0 26 27 0 0 2
1811 508
1621 508
16 12 21 0 0 4224 0 27 26 0 0 2
1621 499
1811 499
15 11 22 0 0 4224 0 27 26 0 0 2
1621 490
1811 490
9 0 47 0 0 0 0 26 0 0 110 2
1805 454
1801 454
1 10 47 0 0 0 0 3 26 0 0 3
1801 426
1801 463
1805 463
3 0 2 0 0 0 0 26 0 0 112 3
1881 472
1895 472
1895 463
2 0 2 0 0 0 0 26 0 0 113 3
1881 463
1903 463
1903 456
1 1 2 0 0 0 0 26 19 0 0 3
1875 454
1875 456
1922 456
1 8 48 0 0 8320 0 25 26 0 0 3
2096 455
2096 517
1875 517
2 7 49 0 0 8320 0 25 26 0 0 3
2090 455
2090 508
1875 508
3 6 50 0 0 8320 0 25 26 0 0 3
2084 455
2084 499
1875 499
4 5 51 0 0 8320 0 25 26 0 0 3
2078 455
2078 490
1875 490
2 4 52 0 0 12416 0 24 26 0 0 4
1965 464
1954 464
1954 481
1875 481
8 1 53 0 0 8320 0 25 24 0 0 3
2054 455
2054 464
1995 464
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1759 368 1871 389
1768 375 1872 390
13 Write control
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1160 565 1192 586
1168 572 1192 587
3 SW2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1308 592 1340 613
1317 598 1341 613
3 SW3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1356 403 1388 424
1364 410 1388 425
3 SW1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1793 377 1825 398
1802 383 1826 398
3 SW4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1328 388 1440 409
1337 394 1441 409
13 Reset control
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
1114 597 1234 618
1123 603 1235 618
14 pulser control
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1291 610 1403 631
1299 617 1403 632
13 clock control
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
