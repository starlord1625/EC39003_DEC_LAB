CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
530 50 2 100 9
0 71 1536 864
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 864
143654930 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 1395 390 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
2 +V
167 976 80 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 1392 483 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 74LS157
122 1437 426 0 14 29
0 4 7 15 14 14 6 13 5 12
2 8 9 10 11
0
0 0 13040 0
7 74LS157
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
6153 0 0
0
0
10 4-In NAND~
219 1268 546 0 5 22
0 19 18 17 16 5
0
0 0 624 0
6 74LS20
-21 -28 21 -20
3 U6B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 -1768304749
65 0 0 0 2 2 4 0
1 U
5394 0 0
0
0
10 2-In NAND~
219 1265 459 0 3 22
0 18 20 6
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -1650864232
65 0 0 0 4 1 5 0
1 U
7734 0 0
0
0
10 4-In NAND~
219 1246 372 0 5 22
0 22 21 20 16 7
0
0 0 624 0
6 74LS20
-21 -28 21 -20
3 U6A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 -1701195873
65 0 0 0 2 1 4 0
1 U
9914 0 0
0
0
7 Ground~
168 948 664 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
9 Inverter~
13 1148 477 0 2 22
0 18 13
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 3 0
1 U
3549 0 0
0
0
10 3-In NAND~
219 1168 507 0 4 22
0 19 18 17 12
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 2 0
1 U
7931 0 0
0
0
10 3-In NAND~
219 1168 449 0 4 22
0 18 17 20 14
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 2 0
1 U
9325 0 0
0
0
10 3-In NAND~
219 1165 402 0 4 22
0 22 21 16 15
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
8903 0 0
0
0
7 74LS138
19 1002 607 0 14 29
0 24 25 26 36 2 2 16 20 23
21 17 18 19 22
0
0 0 13296 602
7 74LS138
51 -3 100 5
2 U3
69 -13 83 -5
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
7 Pulser~
4 931 785 0 10 12
0 37 38 27 39 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3363 0 0
0
0
6 74LS93
109 1013 703 0 8 17
0 2 2 27 26 40 24 25 26
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U1
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
7 Ground~
168 1017 762 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
9 CA 7-Seg~
184 1021 156 0 18 19
10 29 30 31 32 33 34 35 41 28
2 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3874 0 0
0
0
6 74LS47
187 994 291 0 14 29
0 11 10 9 8 42 43 35 34 33
32 31 30 29 27
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U2
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6671 0 0
0
0
9 Resistor~
219 1021 96 0 4 5
0 28 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
66
1 2 3 0 0 4224 0 2 19 0 0 4
976 89
1004 89
1004 78
1021 78
1 1 4 0 0 4224 0 1 4 0 0 2
1407 390
1405 390
5 8 5 0 0 8320 0 5 4 0 0 4
1295 546
1355 546
1355 453
1405 453
3 6 6 0 0 8320 0 6 4 0 0 3
1292 459
1292 435
1405 435
5 2 7 0 0 4224 0 7 4 0 0 4
1273 372
1357 372
1357 399
1405 399
10 1 2 0 0 4096 0 4 3 0 0 4
1399 471
1390 471
1390 477
1392 477
4 11 8 0 0 16512 0 18 4 0 0 7
1008 328
1008 348
1168 348
1168 332
1486 332
1486 408
1469 408
3 12 9 0 0 16512 0 18 4 0 0 7
1017 328
1017 345
1151 345
1151 320
1502 320
1502 426
1469 426
2 13 10 0 0 16512 0 18 4 0 0 7
1026 328
1026 341
1144 341
1144 309
1519 309
1519 444
1469 444
1 14 11 0 0 12416 0 18 4 0 0 6
1035 328
1128 328
1128 298
1540 298
1540 462
1469 462
4 9 12 0 0 4224 0 10 4 0 0 4
1195 507
1340 507
1340 462
1405 462
2 7 13 0 0 12416 0 9 4 0 0 6
1169 477
1212 477
1212 493
1315 493
1315 444
1405 444
0 5 14 0 0 8192 0 0 4 14 0 3
1389 417
1389 426
1405 426
4 4 14 0 0 8320 0 11 4 0 0 3
1195 449
1195 417
1405 417
4 3 15 0 0 4224 0 12 4 0 0 4
1192 402
1353 402
1353 408
1405 408
4 0 16 0 0 4224 0 5 0 0 43 2
1244 560
1026 560
3 0 17 0 0 4224 0 5 0 0 47 2
1244 551
990 551
2 0 18 0 0 4224 0 5 0 0 48 2
1244 542
981 542
1 0 19 0 0 4224 0 5 0 0 49 2
1244 533
972 533
0 1 18 0 0 0 0 0 6 28 0 5
1109 477
1109 466
1233 466
1233 450
1241 450
0 2 20 0 0 4224 0 0 6 44 0 3
1017 486
1241 486
1241 468
4 0 16 0 0 0 0 7 0 0 43 2
1222 386
1026 386
0 3 20 0 0 0 0 0 7 44 0 4
1017 373
1215 373
1215 377
1222 377
0 2 21 0 0 8320 0 0 7 46 0 4
999 371
999 363
1222 363
1222 368
1 0 22 0 0 4224 0 7 0 0 50 3
1222 359
963 359
963 367
6 5 2 0 0 0 0 13 13 0 0 2
963 642
972 642
6 1 2 0 0 8192 0 13 8 0 0 3
963 642
948 642
948 658
0 1 18 0 0 0 0 0 9 48 0 3
981 478
981 477
1133 477
2 0 18 0 0 0 0 10 0 0 35 2
1144 507
1144 507
2 0 17 0 0 0 0 11 0 0 39 2
1144 449
1144 448
3 0 16 0 0 0 0 12 0 0 40 2
1141 411
1141 411
2 0 21 0 0 0 0 12 0 0 41 2
1141 402
1141 402
1 0 22 0 0 0 0 12 0 0 42 2
1141 393
1141 393
3 0 17 0 0 0 0 10 0 0 47 2
1144 516
990 516
0 0 18 0 0 0 0 0 0 0 48 2
1148 507
981 507
1 0 19 0 0 0 0 10 0 0 49 2
1144 498
972 498
1 0 18 0 0 0 0 11 0 0 48 3
1144 440
1144 439
981 439
3 0 20 0 0 0 0 11 0 0 44 3
1144 458
1144 457
1017 457
0 0 17 0 0 0 0 0 0 0 47 2
1148 448
990 448
0 0 16 0 0 0 0 0 0 0 43 2
1145 411
1026 411
0 0 21 0 0 0 0 0 0 0 46 2
1146 402
999 402
0 0 22 0 0 0 0 0 0 0 50 2
1145 393
963 393
7 0 16 0 0 0 0 13 0 0 0 2
1026 566
1026 366
8 0 20 0 0 0 0 13 0 0 0 2
1017 566
1017 364
9 0 23 0 0 4224 0 13 0 0 0 2
1008 566
1008 372
10 0 21 0 0 0 0 13 0 0 0 2
999 566
999 368
11 0 17 0 0 0 0 13 0 0 0 2
990 566
990 365
12 0 18 0 0 0 0 13 0 0 0 2
981 566
981 361
13 0 19 0 0 0 0 13 0 0 0 2
972 566
972 366
14 0 22 0 0 0 0 13 0 0 0 2
963 566
963 363
6 1 24 0 0 12416 0 15 13 0 0 4
1011 669
1011 653
1026 653
1026 636
7 2 25 0 0 4224 0 15 13 0 0 4
1002 669
1002 643
1017 643
1017 636
0 3 26 0 0 4096 0 0 13 55 0 3
993 662
993 636
1008 636
14 0 27 0 0 12416 0 18 0 0 56 6
954 264
954 236
712 236
712 740
963 740
963 776
4 8 26 0 0 12416 0 15 15 0 0 6
993 739
993 752
970 752
970 662
993 662
993 669
3 3 27 0 0 0 0 15 14 0 0 3
1002 739
1002 776
955 776
1 0 2 0 0 4224 0 15 0 0 58 3
1020 733
1020 752
1015 752
2 1 2 0 0 0 0 15 16 0 0 4
1011 733
1011 752
1017 752
1017 756
9 1 28 0 0 4224 0 17 19 0 0 2
1021 120
1021 114
13 1 29 0 0 12416 0 18 17 0 0 5
981 258
981 227
1001 227
1001 192
1000 192
12 2 30 0 0 12416 0 18 17 0 0 5
990 258
990 235
1007 235
1007 192
1006 192
11 3 31 0 0 12416 0 18 17 0 0 5
999 258
999 245
1013 245
1013 192
1012 192
4 10 32 0 0 16512 0 17 18 0 0 7
1018 192
1019 192
1019 196
1017 196
1017 251
1008 251
1008 258
5 9 33 0 0 16512 0 17 18 0 0 6
1024 192
1025 192
1025 199
1021 199
1021 258
1017 258
8 6 34 0 0 4224 0 18 17 0 0 5
1026 258
1026 203
1031 203
1031 192
1030 192
7 7 35 0 0 12416 0 17 18 0 0 4
1036 192
1036 190
1035 190
1035 258
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
