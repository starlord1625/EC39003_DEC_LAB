CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1070 30 5 120 9
0 71 1536 864
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 864
143654930 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 1789 426 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 1326 584 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 1183 557 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 1369 453 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
7 Ground~
168 1521 442 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 1652 431 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 1922 462 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
8 2-In OR~
219 1368 532 0 3 22
0 6 7 3
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1330618039
65 0 0 0 4 1 3 0
1 U
3747 0 0
0
0
7 Pulser~
4 1200 502 0 10 12
0 32 33 4 34 0 0 5 5 3
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3549 0 0
0
0
9 2-In AND~
219 1280 530 0 3 22
0 4 5 6
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
7931 0 0
0
0
6 74LS93
109 1462 507 0 8 17
0 8 8 35 3 11 10 9 36
0
0 0 13024 0
6 74LS93
-21 -35 21 -27
2 U5
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
7 Buffer~
58 1980 464 0 2 22
0 22 21
0
0 0 608 180
4 4050
-14 -19 14 -11
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
8903 0 0
0
0
10 Ascii Key~
169 2075 431 0 11 12
0 17 18 19 20 37 38 39 22 0
0 49
0
0 0 4640 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3834 0 0
0
0
7 74LS173
129 1843 481 0 14 29
0 2 2 2 21 20 19 18 17 12
12 14 13 15 16
0
0 0 13024 512
7 74LS173
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
6 1K RAM
79 1589 472 0 20 41
0 2 2 2 2 2 2 2 11 10
9 40 41 42 43 14 13 15 16 2
12
0
0 0 13024 0
5 RAM1K
-17 -19 18 -11
2 U1
-7 -70 7 -62
0
15 DVCC=22;DGND=11
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
6 74LS47
187 1700 317 0 14 29
0 14 13 15 16 44 45 31 30 29
28 27 26 25 3
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
2 U2
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4718 0 0
0
0
9 CA 7-Seg~
184 1727 182 0 18 19
10 25 26 27 28 29 30 31 46 24
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3874 0 0
0
0
2 +V
167 1727 72 0 1 3
0 23
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6671 0 0
0
0
9 Resistor~
219 1727 122 0 4 5
0 24 23 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
48
0 14 3 0 0 4224 0 0 16 6 0 4
1407 532
1407 279
1660 279
1660 290
3 1 4 0 0 8320 0 9 10 0 0 4
1224 493
1238 493
1238 521
1256 521
1 2 5 0 0 4224 0 3 10 0 0 4
1195 557
1238 557
1238 539
1256 539
3 1 6 0 0 8320 0 10 8 0 0 3
1301 530
1301 523
1355 523
2 1 7 0 0 8320 0 8 2 0 0 4
1355 541
1345 541
1345 584
1338 584
3 4 3 0 0 0 0 8 11 0 0 3
1401 532
1424 532
1424 525
0 1 8 0 0 8192 0 0 11 8 0 3
1415 497
1415 498
1430 498
1 2 8 0 0 8320 0 4 11 0 0 4
1381 453
1415 453
1415 507
1430 507
7 10 9 0 0 8320 0 11 15 0 0 3
1494 516
1494 517
1557 517
6 9 10 0 0 8320 0 11 15 0 0 3
1494 507
1494 508
1557 508
8 5 11 0 0 8320 0 15 11 0 0 3
1557 499
1557 498
1494 498
2 0 2 0 0 4096 0 15 0 0 17 2
1557 445
1532 445
3 0 2 0 0 0 0 15 0 0 17 2
1557 454
1532 454
4 0 2 0 0 0 0 15 0 0 17 2
1557 463
1532 463
5 0 2 0 0 0 0 15 0 0 17 2
1557 472
1532 472
6 0 2 0 0 0 0 15 0 0 17 2
1557 481
1532 481
0 7 2 0 0 4224 0 0 15 18 0 3
1532 436
1532 490
1557 490
1 1 2 0 0 0 0 5 15 0 0 2
1521 436
1557 436
19 1 2 0 0 0 0 15 6 0 0 4
1627 436
1627 420
1652 420
1652 425
20 0 12 0 0 4224 0 15 0 0 30 2
1627 445
1801 445
2 0 13 0 0 4096 0 16 0 0 27 2
1732 354
1732 499
1 0 14 0 0 4096 0 16 0 0 28 2
1741 354
1741 490
3 0 15 0 0 4096 0 16 0 0 26 2
1723 354
1723 508
4 0 16 0 0 4096 0 16 0 0 25 2
1714 354
1714 517
18 14 16 0 0 4224 0 15 14 0 0 2
1621 517
1811 517
13 17 15 0 0 4224 0 14 15 0 0 2
1811 508
1621 508
16 12 13 0 0 4224 0 15 14 0 0 2
1621 499
1811 499
15 11 14 0 0 4224 0 15 14 0 0 2
1621 490
1811 490
9 0 12 0 0 0 0 14 0 0 30 2
1805 454
1801 454
1 10 12 0 0 0 0 1 14 0 0 3
1801 426
1801 463
1805 463
3 0 2 0 0 0 0 14 0 0 32 3
1881 472
1895 472
1895 463
2 0 2 0 0 0 0 14 0 0 33 3
1881 463
1903 463
1903 456
1 1 2 0 0 0 0 14 7 0 0 3
1875 454
1875 456
1922 456
1 8 17 0 0 8320 0 13 14 0 0 3
2096 455
2096 517
1875 517
2 7 18 0 0 8320 0 13 14 0 0 3
2090 455
2090 508
1875 508
3 6 19 0 0 8320 0 13 14 0 0 3
2084 455
2084 499
1875 499
4 5 20 0 0 8320 0 13 14 0 0 3
2078 455
2078 490
1875 490
2 4 21 0 0 12416 0 12 14 0 0 4
1965 464
1954 464
1954 481
1875 481
8 1 22 0 0 8320 0 13 12 0 0 3
2054 455
2054 464
1995 464
1 2 23 0 0 4224 0 18 19 0 0 2
1727 81
1727 104
9 1 24 0 0 4224 0 17 19 0 0 2
1727 146
1727 140
13 1 25 0 0 12416 0 16 17 0 0 5
1687 284
1687 253
1707 253
1707 218
1706 218
12 2 26 0 0 12416 0 16 17 0 0 5
1696 284
1696 261
1713 261
1713 218
1712 218
11 3 27 0 0 12416 0 16 17 0 0 5
1705 284
1705 271
1719 271
1719 218
1718 218
4 10 28 0 0 16512 0 17 16 0 0 7
1724 218
1725 218
1725 222
1723 222
1723 277
1714 277
1714 284
5 9 29 0 0 16512 0 17 16 0 0 6
1730 218
1731 218
1731 225
1727 225
1727 284
1723 284
8 6 30 0 0 4224 0 16 17 0 0 5
1732 284
1732 229
1737 229
1737 218
1736 218
7 7 31 0 0 12416 0 17 16 0 0 4
1742 218
1742 216
1741 216
1741 284
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1291 610 1403 631
1299 617 1403 632
13 clock control
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
1114 597 1234 618
1123 603 1235 618
14 pulser control
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1328 388 1440 409
1337 394 1441 409
13 Reset control
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1759 368 1871 389
1768 375 1872 390
13 Write control
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1793 377 1825 398
1802 383 1826 398
3 SW4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1356 403 1388 424
1364 410 1388 425
3 SW1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1308 592 1340 613
1317 598 1341 613
3 SW3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1160 565 1192 586
1168 572 1192 587
3 SW2
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
