CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1000 70 2 80 9
0 76 1536 869
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 76 1536 869
143654930 0
0
6 Title:
5 Name:
0
0
0
32
13 Logic Switch~
5 1705 843 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 1639 809 0 1 11
0 34
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 1557 781 0 1 11
0 33
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V9
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 1504 755 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V8
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 1066 754 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 1061 804 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 1065 857 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 1060 907 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 1115 984 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3549 0 0
0
0
8 3-In OR~
219 1391 538 0 4 22
0 3 5 4 9
0
0 0 624 90
4 4075
-14 -24 14 -16
3 U8A
28 -3 49 5
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
7931 0 0
0
0
9 2-In AND~
219 1416 597 0 3 22
0 7 8 4
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U6D
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 -170575095
65 0 0 0 4 4 3 0
1 U
9325 0 0
0
0
9 2-In AND~
219 1374 599 0 3 22
0 6 8 5
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U6C
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 -120243452
65 0 0 0 4 3 3 0
1 U
8903 0 0
0
0
7 Ground~
168 1543 526 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
7 Ground~
168 1817 659 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
6 74LS83
105 1803 552 0 14 29
0 8 6 7 14 2 15 15 2 2
13 12 11 10 52
0
0 0 13040 90
7 74LS83A
-24 -60 25 -52
2 U9
57 -3 71 5
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
7 Ground~
168 1262 379 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
7 74LS157
122 1593 462 0 14 29
0 9 10 14 11 7 12 6 13 8
2 19 18 17 16
0
0 0 13040 602
7 74LS157
-24 -60 25 -52
2 U7
54 -6 68 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3874 0 0
0
0
9 2-In AND~
219 1339 635 0 3 22
0 21 20 3
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U6A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -120243452
65 0 0 0 4 1 3 0
1 U
6671 0 0
0
0
9 Inverter~
13 1306 681 0 2 22
0 22 21
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 2 0
1 U
3789 0 0
0
0
9 2-In XOR~
219 1190 762 0 3 22
0 26 22 28
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
4871 0 0
0
0
9 2-In XOR~
219 1190 813 0 3 22
0 27 22 29
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 1 0
1 U
3750 0 0
0
0
9 2-In XOR~
219 1188 915 0 3 22
0 25 22 31
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
8778 0 0
0
0
9 2-In XOR~
219 1189 865 0 3 22
0 24 22 30
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -204129521
65 0 0 0 4 1 1 0
1 U
538 0 0
0
0
6 74LS83
105 1412 696 0 14 29
0 32 33 34 23 28 29 30 31 22
8 6 7 14 20
0
0 0 13040 602
7 74LS83A
-24 -60 25 -52
2 U3
57 -3 71 5
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6843 0 0
0
0
2 +V
167 1600 59 0 1 3
0 15
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3136 0 0
0
0
9 CA 7-Seg~
184 1600 169 0 18 19
10 36 37 38 39 40 41 42 53 35
0 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5950 0 0
0
0
6 74LS47
187 1573 304 0 14 29
0 16 17 18 19 54 55 42 41 40
39 38 37 36 56
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
6 74LS47
187 1225 300 0 14 29
0 2 2 2 9 57 58 51 50 49
48 47 46 45 59
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U2
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6828 0 0
0
0
9 CA 7-Seg~
184 1252 165 0 18 19
10 45 46 47 48 49 50 51 60 44
2 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6735 0 0
0
0
2 +V
167 1252 55 0 1 3
0 43
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8365 0 0
0
0
9 Resistor~
219 1600 109 0 4 5
0 35 15 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 1252 105 0 4 5
0 44 43 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
75
3 1 3 0 0 8320 0 18 10 0 0 4
1338 611
1338 567
1385 567
1385 554
3 3 4 0 0 4224 0 10 11 0 0 3
1403 554
1403 573
1415 573
3 2 5 0 0 8320 0 12 10 0 0 3
1373 575
1394 575
1394 553
1 0 6 0 0 8192 0 12 0 0 32 3
1364 620
1364 649
1414 649
1 0 7 0 0 8192 0 11 0 0 33 3
1406 618
1408 618
1408 635
2 0 8 0 0 8192 0 11 0 0 7 3
1424 618
1423 618
1423 656
2 0 8 0 0 8192 0 12 0 0 31 3
1382 620
1382 656
1423 656
10 1 2 0 0 4096 0 17 13 0 0 4
1547 499
1547 514
1543 514
1543 520
4 0 9 0 0 8320 0 28 0 0 30 4
1239 337
1239 459
1417 459
1417 508
2 13 10 0 0 8320 0 17 15 0 0 4
1619 493
1619 503
1819 503
1819 522
4 12 11 0 0 8320 0 17 15 0 0 4
1601 493
1601 510
1810 510
1810 522
6 11 12 0 0 8320 0 17 15 0 0 4
1583 493
1583 517
1801 517
1801 522
8 10 13 0 0 8320 0 17 15 0 0 3
1565 493
1565 522
1792 522
0 1 8 0 0 4224 0 0 15 31 0 3
1553 653
1765 653
1765 586
0 2 6 0 0 4224 0 0 15 32 0 3
1573 644
1774 644
1774 586
0 3 7 0 0 4224 0 0 15 33 0 3
1590 633
1783 633
1783 586
0 4 14 0 0 4096 0 0 15 34 0 3
1609 626
1792 626
1792 586
6 0 15 0 0 4096 0 15 0 0 19 3
1810 586
1810 604
1819 604
0 7 15 0 0 8320 0 0 15 58 0 5
1600 82
2007 82
2007 604
1819 604
1819 586
9 0 2 0 0 4096 0 15 0 0 21 3
1846 586
1846 624
1828 624
8 1 2 0 0 4224 0 15 14 0 0 3
1828 586
1828 653
1817 653
5 1 2 0 0 0 0 15 14 0 0 3
1801 586
1801 653
1817 653
1 0 2 0 0 0 0 28 0 0 24 3
1266 337
1266 359
1257 359
2 0 2 0 0 0 0 28 0 0 25 2
1257 337
1257 373
3 1 2 0 0 0 0 28 16 0 0 3
1248 337
1248 373
1262 373
14 1 16 0 0 8320 0 17 27 0 0 4
1556 429
1556 390
1614 390
1614 341
13 2 17 0 0 12416 0 17 27 0 0 4
1574 429
1574 401
1605 401
1605 341
3 12 18 0 0 4224 0 27 17 0 0 4
1596 341
1596 422
1592 422
1592 429
4 11 19 0 0 4224 0 27 17 0 0 4
1587 341
1587 408
1610 408
1610 429
1 4 9 0 0 0 0 17 10 0 0 5
1628 493
1628 545
1461 545
1461 508
1394 508
10 9 8 0 0 0 0 24 17 0 0 4
1423 666
1423 653
1556 653
1556 493
11 7 6 0 0 0 0 24 17 0 0 4
1414 666
1414 644
1574 644
1574 493
12 5 7 0 0 0 0 24 17 0 0 5
1405 666
1408 666
1408 633
1592 633
1592 493
13 3 14 0 0 8320 0 24 17 0 0 4
1396 666
1396 626
1610 626
1610 493
2 14 20 0 0 8320 0 18 24 0 0 3
1347 656
1347 666
1369 666
2 1 21 0 0 4224 0 19 18 0 0 3
1309 663
1329 663
1329 656
1 0 22 0 0 8192 0 19 0 0 38 3
1309 699
1309 746
1369 746
0 9 22 0 0 4224 0 0 24 49 0 3
1127 966
1369 966
1369 730
1 0 23 0 0 0 0 1 0 0 57 2
1693 843
1693 843
1 0 24 0 0 4096 0 7 0 0 44 2
1077 857
1077 856
1 0 25 0 0 4096 0 8 0 0 45 2
1072 907
1072 906
1 1 26 0 0 4224 0 20 5 0 0 3
1174 753
1078 753
1078 754
1 1 27 0 0 4224 0 21 6 0 0 2
1174 804
1073 804
1 0 24 0 0 4224 0 23 0 0 0 2
1173 856
1072 856
1 0 25 0 0 4224 0 22 0 0 0 2
1172 906
1069 906
0 2 22 0 0 0 0 0 20 47 0 3
1132 823
1132 771
1174 771
0 2 22 0 0 0 0 0 21 48 0 3
1132 874
1132 822
1174 822
0 2 22 0 0 0 0 0 23 49 0 3
1128 924
1128 874
1173 874
2 1 22 0 0 0 0 22 9 0 0 3
1172 924
1127 924
1127 984
3 5 28 0 0 4224 0 20 24 0 0 3
1223 762
1414 762
1414 730
3 6 29 0 0 4224 0 21 24 0 0 3
1223 813
1405 813
1405 730
3 7 30 0 0 4224 0 23 24 0 0 3
1222 865
1396 865
1396 730
3 8 31 0 0 8320 0 22 24 0 0 3
1221 915
1387 915
1387 730
1 1 32 0 0 8320 0 24 4 0 0 4
1450 730
1450 756
1492 756
1492 755
2 1 33 0 0 8320 0 24 3 0 0 3
1441 730
1441 781
1545 781
3 1 34 0 0 8320 0 24 2 0 0 4
1432 730
1432 808
1627 808
1627 809
4 0 23 0 0 8320 0 24 0 0 0 3
1423 730
1423 843
1699 843
1 2 15 0 0 0 0 25 31 0 0 2
1600 68
1600 91
9 1 35 0 0 4224 0 26 31 0 0 2
1600 133
1600 127
13 1 36 0 0 12416 0 27 26 0 0 5
1560 271
1560 240
1580 240
1580 205
1579 205
12 2 37 0 0 12416 0 27 26 0 0 5
1569 271
1569 248
1586 248
1586 205
1585 205
11 3 38 0 0 12416 0 27 26 0 0 5
1578 271
1578 258
1592 258
1592 205
1591 205
4 10 39 0 0 16512 0 26 27 0 0 7
1597 205
1598 205
1598 209
1596 209
1596 264
1587 264
1587 271
5 9 40 0 0 16512 0 26 27 0 0 6
1603 205
1604 205
1604 212
1600 212
1600 271
1596 271
8 6 41 0 0 4224 0 27 26 0 0 5
1605 271
1605 216
1610 216
1610 205
1609 205
7 7 42 0 0 12416 0 26 27 0 0 4
1615 205
1615 203
1614 203
1614 271
1 2 43 0 0 4224 0 30 32 0 0 2
1252 64
1252 87
9 1 44 0 0 4224 0 29 32 0 0 2
1252 129
1252 123
13 1 45 0 0 12416 0 28 29 0 0 5
1212 267
1212 236
1232 236
1232 201
1231 201
12 2 46 0 0 12416 0 28 29 0 0 5
1221 267
1221 244
1238 244
1238 201
1237 201
11 3 47 0 0 12416 0 28 29 0 0 5
1230 267
1230 254
1244 254
1244 201
1243 201
4 10 48 0 0 16512 0 29 28 0 0 7
1249 201
1250 201
1250 205
1248 205
1248 260
1239 260
1239 267
5 9 49 0 0 16512 0 29 28 0 0 6
1255 201
1256 201
1256 208
1252 208
1252 267
1248 267
8 6 50 0 0 4224 0 28 29 0 0 5
1257 267
1257 212
1262 212
1262 201
1261 201
7 7 51 0 0 12416 0 29 28 0 0 4
1267 201
1267 199
1266 199
1266 267
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
