CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
600 110 3 120 9
0 71 1536 864
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 864
177209362 0
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 983 362 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 1003 323 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 1269 564 0 10 11
0 41 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
7 Ground~
168 1013 244 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
10 Ascii Key~
169 906 247 0 11 12
0 6 5 4 3 43 44 45 46 0
0 57
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
5394 0 0
0
0
9 Inverter~
13 1125 540 0 2 22
0 17 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 3 0
1 U
7734 0 0
0
0
6 74LS95
110 1088 303 0 12 25
0 18 17 17 6 5 4 3 2 7
47 48 49
0
0 0 13040 692
6 74LS95
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
9914 0 0
0
0
9 2-In AND~
219 1442 329 0 3 22
0 26 7 19
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
3747 0 0
0
0
9 2-In AND~
219 1388 330 0 3 22
0 25 7 20
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
3549 0 0
0
0
9 2-In AND~
219 1340 330 0 3 22
0 24 7 21
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
7931 0 0
0
0
9 2-In AND~
219 1288 327 0 3 22
0 23 7 22
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1612193530
65 0 0 0 4 1 2 0
1 U
9325 0 0
0
0
7 74LS173
129 1547 221 0 14 29
0 2 2 2 31 30 29 28 27 2
2 23 24 25 26
0
0 0 13040 512
7 74LS173
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
10 Ascii Key~
169 1779 171 0 11 12
0 27 28 29 30 50 51 52 32 0
0 56
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3834 0 0
0
0
7 Buffer~
58 1684 204 0 2 22
0 32 31
0
0 0 624 180
4 4050
-14 -19 14 -11
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
3363 0 0
0
0
7 Ground~
168 1626 202 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
7 Ground~
168 1490 176 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
14 Logic Display~
6 1194 696 0 1 2
10 35
0
0 0 53872 180
6 100MEG
3 -16 45 -8
4 W128
5 0 33 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 1258 698 0 1 2
10 33
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 W64
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 1315 701 0 1 2
10 36
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 W32
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 1368 702 0 1 2
10 37
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 W16
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 1422 704 0 1 2
10 38
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 W8
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3750 0 0
0
0
14 Logic Display~
6 1471 704 0 1 2
10 39
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 W4
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8778 0 0
0
0
14 Logic Display~
6 1519 705 0 1 2
10 40
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 W2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
538 0 0
0
0
14 Logic Display~
6 1564 707 0 1 2
10 34
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 W1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6843 0 0
0
0
7 Ground~
168 1399 430 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3136 0 0
0
0
7 74LS273
150 1355 591 0 18 37
0 41 16 8 9 10 11 12 13 14
15 35 33 36 37 38 39 40 34
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
2 U9
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
5950 0 0
0
0
6 74LS83
105 1462 480 0 14 29
0 38 39 40 34 2 2 2 2 2
13 14 15 53 42
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U8
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
6 74LS83
105 1285 475 0 14 29
0 35 33 36 37 22 21 20 19 42
9 10 11 12 8
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U5
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6828 0 0
0
0
64
4 7 3 0 0 8320 0 5 7 0 0 3
909 271
909 280
1056 280
3 6 4 0 0 8320 0 5 7 0 0 3
915 271
915 289
1056 289
2 5 5 0 0 8320 0 5 7 0 0 3
921 271
921 298
1056 298
1 4 6 0 0 8320 0 5 7 0 0 3
927 271
927 307
1056 307
2 0 7 0 0 4096 0 9 0 0 8 2
1377 308
1377 288
0 0 7 0 0 4096 0 0 0 8 7 3
1329 291
1274 291
1274 298
9 2 7 0 0 4224 0 7 11 0 0 3
1120 298
1277 298
1277 305
2 2 7 0 0 0 0 8 10 0 0 4
1431 307
1431 288
1329 288
1329 308
8 1 2 0 0 8192 0 7 4 0 0 5
1056 271
1036 271
1036 234
1013 234
1013 238
14 3 8 0 0 4224 0 28 26 0 0 4
1328 509
1328 558
1332 558
1332 564
10 4 9 0 0 8320 0 28 26 0 0 4
1274 509
1274 543
1341 543
1341 564
11 5 10 0 0 8320 0 28 26 0 0 4
1283 509
1283 535
1350 535
1350 564
12 6 11 0 0 8320 0 28 26 0 0 4
1292 509
1292 529
1359 529
1359 564
13 7 12 0 0 8320 0 28 26 0 0 4
1301 509
1301 523
1368 523
1368 564
10 8 13 0 0 8320 0 27 26 0 0 4
1473 514
1473 548
1377 548
1377 564
9 11 14 0 0 8320 0 26 27 0 0 4
1386 564
1386 553
1464 553
1464 514
12 10 15 0 0 8320 0 27 26 0 0 3
1455 514
1455 564
1395 564
2 2 16 0 0 4224 0 6 26 0 0 5
1146 540
1249 540
1249 548
1323 548
1323 564
0 1 17 0 0 4224 0 0 6 22 0 3
1028 325
1028 540
1110 540
1 1 18 0 0 4224 0 1 7 0 0 3
995 362
1056 362
1056 334
3 0 17 0 0 0 0 7 0 0 22 3
1050 316
1035 316
1035 325
1 2 17 0 0 0 0 2 7 0 0 3
1015 323
1015 325
1050 325
5 0 2 0 0 8192 0 27 0 0 54 3
1464 450
1464 424
1419 424
6 0 2 0 0 0 0 27 0 0 54 3
1455 450
1455 431
1419 431
7 0 2 0 0 0 0 27 0 0 54 3
1446 450
1446 440
1419 440
8 0 2 0 0 0 0 27 0 0 54 3
1437 450
1437 445
1419 445
8 3 19 0 0 8320 0 28 8 0 0 6
1310 445
1310 401
1396 401
1396 362
1440 362
1440 352
7 3 20 0 0 8320 0 28 9 0 0 4
1301 445
1301 387
1386 387
1386 353
6 3 21 0 0 4224 0 28 10 0 0 4
1292 445
1292 374
1338 374
1338 353
3 5 22 0 0 8320 0 11 28 0 0 3
1286 350
1283 350
1283 445
11 1 23 0 0 4224 0 12 11 0 0 3
1515 230
1295 230
1295 305
12 1 24 0 0 4224 0 12 10 0 0 3
1515 239
1347 239
1347 308
13 1 25 0 0 4224 0 12 9 0 0 3
1515 248
1395 248
1395 308
14 1 26 0 0 4224 0 12 8 0 0 3
1515 257
1449 257
1449 307
9 0 2 0 0 0 0 12 0 0 36 2
1509 194
1505 194
1 10 2 0 0 0 0 16 12 0 0 5
1490 170
1490 166
1505 166
1505 203
1509 203
3 0 2 0 0 0 0 12 0 0 38 3
1585 212
1599 212
1599 203
2 0 2 0 0 0 0 12 0 0 39 3
1585 203
1607 203
1607 196
1 1 2 0 0 8320 0 12 15 0 0 3
1579 194
1579 196
1626 196
1 8 27 0 0 8320 0 13 12 0 0 3
1800 195
1800 257
1579 257
2 7 28 0 0 8320 0 13 12 0 0 3
1794 195
1794 248
1579 248
3 6 29 0 0 8320 0 13 12 0 0 3
1788 195
1788 239
1579 239
4 5 30 0 0 8320 0 13 12 0 0 3
1782 195
1782 230
1579 230
2 4 31 0 0 12416 0 14 12 0 0 4
1669 204
1658 204
1658 221
1579 221
8 1 32 0 0 8320 0 13 14 0 0 3
1758 195
1758 204
1699 204
1 0 33 0 0 4096 0 18 0 0 58 2
1258 684
1258 640
0 1 34 0 0 4096 0 0 24 63 0 4
1532 628
1532 683
1564 683
1564 693
0 1 35 0 0 4096 0 0 17 59 0 3
1233 631
1233 682
1194 682
0 1 36 0 0 8192 0 0 19 57 0 3
1313 651
1315 651
1315 687
0 1 37 0 0 4096 0 0 20 56 0 3
1356 662
1356 688
1368 688
1 0 38 0 0 4096 0 21 0 0 60 2
1422 690
1422 662
1 0 39 0 0 4096 0 22 0 0 61 2
1471 690
1471 653
0 1 40 0 0 4096 0 0 23 62 0 2
1519 644
1519 691
1 9 2 0 0 0 0 25 27 0 0 3
1399 424
1419 424
1419 450
1 1 41 0 0 4224 0 26 3 0 0 3
1314 558
1281 558
1281 564
4 14 37 0 0 12416 0 28 26 0 0 6
1274 445
1274 413
1186 413
1186 662
1359 662
1359 628
3 13 36 0 0 12416 0 28 26 0 0 6
1265 445
1265 425
1200 425
1200 651
1350 651
1350 628
2 12 33 0 0 12416 0 28 26 0 0 6
1256 445
1256 438
1219 438
1219 640
1341 640
1341 628
1 11 35 0 0 8320 0 28 26 0 0 5
1247 445
1228 445
1228 631
1332 631
1332 628
15 1 38 0 0 12416 0 26 27 0 0 6
1368 628
1368 662
1585 662
1585 443
1500 443
1500 450
16 2 39 0 0 12416 0 26 27 0 0 6
1377 628
1377 653
1573 653
1573 419
1491 419
1491 450
17 3 40 0 0 12416 0 26 27 0 0 6
1386 628
1386 644
1555 644
1555 428
1482 428
1482 450
18 4 34 0 0 8320 0 26 27 0 0 5
1395 628
1537 628
1537 437
1473 437
1473 450
9 14 42 0 0 8320 0 28 27 0 0 4
1328 445
1386 445
1386 514
1419 514
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1057 545 1129 566
1065 552 1129 567
8 Inverter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
857 352 961 373
865 359 961 374
12 mode control
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
883 307 987 328
891 314 987 329
12 Manual clock
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
868 195 956 216
877 202 957 217
10 Multiplier
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
1730 113 1809 132
1738 119 1810 132
12 Multiplicand
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
1214 566 1299 585
1222 573 1300 586
13 Reset control
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
1598 695 1623 714
1606 702 1624 715
3 LSB
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
1138 690 1163 709
1146 697 1164 710
3 MSB
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 11
1406 601 1479 620
1413 608 1479 621
11 Accumulator
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
