CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
540 150 3 120 9
0 71 1536 864
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 864
177209362 0
0
6 Title:
5 Name:
0
0
0
31
13 Logic Switch~
5 1269 564 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 1022 257 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 901 398 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 804 371 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 1461 263 0 1 11
0 42
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5394 0 0
0
0
14 Logic Display~
6 1194 696 0 1 2
10 4
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L8
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 1258 698 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L7
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 1315 701 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L6
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 1368 702 0 1 2
10 6
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L5
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 1422 704 0 1 2
10 7
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L4
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 1471 704 0 1 2
10 8
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 1519 705 0 1 2
10 9
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 1564 707 0 1 2
10 3
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
7 Ground~
168 1399 430 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3363 0 0
0
0
2 +V
167 1039 199 0 1 3
0 16
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7668 0 0
0
0
7 Ground~
168 1011 316 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4718 0 0
0
0
10 Ascii Key~
169 997 397 0 11 12
0 14 13 12 11 49 50 51 52 0
0 55
0
0 0 4656 0
0
4 KBD2
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3874 0 0
0
0
8 4-In OR~
219 941 491 0 5 22
0 19 20 21 22 18
0
0 0 624 512
4 4072
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0
65 0 0 0 2 1 4 0
1 U
6671 0 0
0
0
7 74LS193
137 1082 378 0 14 29
0 16 10 17 2 11 12 13 14 53
54 22 21 20 19
0
0 0 13040 0
7 74LS193
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3789 0 0
0
0
8 2-In OR~
219 943 346 0 3 22
0 23 24 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 3 0
1 U
4871 0 0
0
0
9 2-In AND~
219 864 331 0 3 22
0 26 25 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3750 0 0
0
0
7 Pulser~
4 674 295 0 10 12
0 55 56 27 57 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8778 0 0
0
0
9 2-In AND~
219 754 323 0 3 22
0 27 18 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
538 0 0
0
0
7 74LS273
150 1355 591 0 18 37
0 15 10 33 34 35 36 29 30 31
32 4 28 5 6 7 8 9 3
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
2 U9
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
6843 0 0
0
0
6 74LS83
105 1462 480 0 14 29
0 7 8 9 3 40 39 38 37 2
29 30 31 32 41
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U8
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3136 0 0
0
0
7 Ground~
168 1341 423 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5950 0 0
0
0
6 74LS83
105 1290 480 0 14 29
0 4 28 5 6 2 2 2 2 41
33 34 35 36 58
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U5
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
7 Ground~
168 1594 299 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6828 0 0
0
0
7 Buffer~
58 1652 301 0 2 22
0 48 47
0
0 0 624 180
4 4050
-14 -19 14 -11
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
6735 0 0
0
0
10 Ascii Key~
169 1747 268 0 11 12
0 43 44 45 46 59 60 61 48 0
0 55
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
8365 0 0
0
0
7 74LS173
129 1515 318 0 14 29
0 2 2 2 47 46 45 44 43 42
42 40 39 38 37
0
0 0 13040 512
7 74LS173
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
4132 0 0
0
0
65
1 0 0 0 0 0 0 7 0 0 32 2
1258 684
1258 640
0 1 3 0 0 4096 0 0 13 37 0 4
1532 628
1532 683
1564 683
1564 693
0 1 4 0 0 4096 0 0 6 33 0 3
1233 631
1233 682
1194 682
0 1 5 0 0 8192 0 0 8 31 0 3
1313 651
1315 651
1315 687
0 1 6 0 0 4096 0 0 9 30 0 3
1356 662
1356 688
1368 688
1 0 7 0 0 4096 0 10 0 0 34 2
1422 690
1422 662
1 0 8 0 0 4096 0 11 0 0 35 2
1471 690
1471 653
0 1 9 0 0 4096 0 0 12 36 0 2
1519 644
1519 691
1 9 2 0 0 8192 0 14 25 0 0 3
1399 424
1419 424
1419 450
0 2 10 0 0 12416 0 0 24 24 0 6
1038 360
1038 297
1166 297
1166 545
1323 545
1323 564
4 5 11 0 0 12416 0 17 19 0 0 5
1000 421
1000 451
1036 451
1036 387
1050 387
3 6 12 0 0 12416 0 17 19 0 0 5
1006 421
1006 439
1042 439
1042 396
1050 396
2 7 13 0 0 8320 0 17 19 0 0 5
1012 421
1012 428
1046 428
1046 405
1050 405
1 8 14 0 0 4224 0 17 19 0 0 3
1018 421
1050 421
1050 414
1 1 15 0 0 4224 0 24 1 0 0 3
1314 558
1281 558
1281 564
1 1 16 0 0 12416 0 15 19 0 0 4
1039 208
1039 206
1050 206
1050 351
1 3 17 0 0 8320 0 2 19 0 0 3
1034 257
1044 257
1044 369
1 4 2 0 0 8320 0 16 19 0 0 4
1011 310
1031 310
1031 378
1050 378
2 5 18 0 0 12416 0 23 18 0 0 4
730 332
718 332
718 491
914 491
1 14 19 0 0 4224 0 18 19 0 0 3
964 478
1114 478
1114 414
13 2 20 0 0 12416 0 19 18 0 0 4
1114 405
1132 405
1132 487
964 487
3 12 21 0 0 4224 0 18 19 0 0 4
964 496
1142 496
1142 396
1114 396
11 4 22 0 0 12416 0 19 18 0 0 4
1114 387
1147 387
1147 505
964 505
3 2 10 0 0 128 0 20 19 0 0 4
976 346
1034 346
1034 360
1050 360
3 1 23 0 0 4224 0 21 20 0 0 4
885 331
920 331
920 337
930 337
2 1 24 0 0 8320 0 20 3 0 0 4
930 355
920 355
920 398
913 398
2 1 25 0 0 8320 0 21 4 0 0 4
840 340
827 340
827 371
816 371
3 1 26 0 0 8320 0 23 21 0 0 3
775 323
775 322
840 322
3 1 27 0 0 8320 0 22 23 0 0 4
698 286
712 286
712 314
730 314
4 14 6 0 0 12416 0 27 24 0 0 6
1279 450
1279 413
1186 413
1186 662
1359 662
1359 628
3 13 5 0 0 12416 0 27 24 0 0 6
1270 450
1270 425
1200 425
1200 651
1350 651
1350 628
2 12 28 0 0 12416 0 27 24 0 0 6
1261 450
1261 438
1219 438
1219 640
1341 640
1341 628
1 11 4 0 0 8320 0 27 24 0 0 5
1252 450
1228 450
1228 631
1332 631
1332 628
15 1 7 0 0 12416 0 24 25 0 0 6
1368 628
1368 662
1585 662
1585 443
1500 443
1500 450
16 2 8 0 0 12416 0 24 25 0 0 6
1377 628
1377 653
1573 653
1573 419
1491 419
1491 450
17 3 9 0 0 12416 0 24 25 0 0 6
1386 628
1386 644
1555 644
1555 428
1482 428
1482 450
18 4 3 0 0 8320 0 24 25 0 0 5
1395 628
1537 628
1537 437
1473 437
1473 450
7 10 29 0 0 8320 0 24 25 0 0 4
1368 564
1368 558
1473 558
1473 514
8 11 30 0 0 8320 0 24 25 0 0 4
1377 564
1377 547
1464 547
1464 514
9 12 31 0 0 8320 0 24 25 0 0 4
1386 564
1386 535
1455 535
1455 514
10 13 32 0 0 8320 0 24 25 0 0 4
1395 564
1395 523
1446 523
1446 514
10 3 33 0 0 8320 0 27 24 0 0 4
1279 514
1279 532
1332 532
1332 564
11 4 34 0 0 8320 0 27 24 0 0 4
1288 514
1288 526
1341 526
1341 564
12 5 35 0 0 8320 0 27 24 0 0 4
1297 514
1297 520
1350 520
1350 564
13 6 36 0 0 4224 0 27 24 0 0 3
1306 514
1359 514
1359 564
8 14 37 0 0 4224 0 25 31 0 0 3
1437 450
1437 354
1483 354
13 7 38 0 0 8320 0 31 25 0 0 3
1483 345
1446 345
1446 450
6 12 39 0 0 4224 0 25 31 0 0 3
1455 450
1455 336
1483 336
11 5 40 0 0 8320 0 31 25 0 0 3
1483 327
1464 327
1464 450
9 14 41 0 0 8320 0 27 25 0 0 4
1333 450
1386 450
1386 514
1419 514
8 0 2 0 0 0 0 27 0 0 54 2
1315 450
1315 408
7 0 2 0 0 0 0 27 0 0 54 2
1306 450
1306 408
6 0 2 0 0 0 0 27 0 0 54 2
1297 450
1297 408
5 1 2 0 0 0 0 27 26 0 0 4
1288 450
1288 408
1341 408
1341 417
9 0 42 0 0 4096 0 31 0 0 56 2
1477 291
1473 291
1 10 42 0 0 4224 0 5 31 0 0 3
1473 263
1473 300
1477 300
3 0 2 0 0 0 0 31 0 0 58 3
1553 309
1567 309
1567 300
2 0 2 0 0 0 0 31 0 0 59 3
1553 300
1575 300
1575 293
1 1 2 0 0 0 0 31 28 0 0 3
1547 291
1547 293
1594 293
1 8 43 0 0 8320 0 30 31 0 0 3
1768 292
1768 354
1547 354
2 7 44 0 0 8320 0 30 31 0 0 3
1762 292
1762 345
1547 345
3 6 45 0 0 8320 0 30 31 0 0 3
1756 292
1756 336
1547 336
4 5 46 0 0 8320 0 30 31 0 0 3
1750 292
1750 327
1547 327
2 4 47 0 0 12416 0 29 31 0 0 4
1637 301
1626 301
1626 318
1547 318
8 1 48 0 0 8320 0 30 29 0 0 3
1726 292
1726 301
1667 301
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
883 406 915 427
892 412 916 427
3 SW3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
859 423 971 444
867 430 971 445
13 clock control
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
634 358 666 379
642 365 666 380
3 SW2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
588 390 708 411
597 396 709 411
14 pulser control
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1465 214 1497 235
1474 220 1498 235
3 SW4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1416 201 1528 222
1424 208 1528 223
13 Write control
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
